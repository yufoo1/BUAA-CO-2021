module CU(
  input  [31:0] io_instr,
  input         io_IsEq,
  output [3:0]  io_ALUOp,
  output        io_WEGRF,
  output        io_WEDM,
  output        io_IsBranchType,
  output        io_IsJType,
  output        io_IsJr,
  output        io_ALUSrc,
  output [1:0]  io_WhichToReg,
  output [1:0]  io_RegDst,
  output        io_IsSignExt
);
  wire [5:0] op = io_instr[31:26]; // @[CU.scala 20:28]
  wire [5:0] func = io_instr[5:0]; // @[CU.scala 21:30]
  wire  RType = op == 6'h0; // @[CU.scala 26:14]
  wire  addu = RType & func == 6'h21; // @[CU.scala 32:25]
  wire  subu = RType & func == 6'h23; // @[CU.scala 38:25]
  wire  ori = op == 6'hd; // @[CU.scala 44:14]
  wire  lw = op == 6'h23; // @[CU.scala 50:14]
  wire  sw = op == 6'h2b; // @[CU.scala 56:14]
  wire  beq = op == 6'h4; // @[CU.scala 62:14]
  wire  lui = op == 6'hf; // @[CU.scala 68:14]
  wire  j = op == 6'h2; // @[CU.scala 74:14]
  wire  jal = op == 6'h3; // @[CU.scala 80:14]
  wire [2:0] _GEN_11 = lui ? 3'h4 : 3'h0; // @[CU.scala 96:31 97:18 99:18]
  wire [2:0] _GEN_12 = ori ? 3'h3 : _GEN_11; // @[CU.scala 94:31 95:18]
  wire [2:0] _GEN_13 = subu ? 3'h1 : _GEN_12; // @[CU.scala 92:25 93:18]
  wire  _T_33 = ori | lui | lw; // @[CU.scala 132:22]
  wire [1:0] _GEN_20 = jal ? 2'h2 : 2'h0; // @[CU.scala 140:31 141:23 143:23]
  assign io_ALUOp = {{1'd0}, _GEN_13};
  assign io_WEGRF = addu | subu | ori | lw | lui | jal; // @[CU.scala 102:41]
  assign io_WEDM = op == 6'h2b; // @[CU.scala 56:14]
  assign io_IsBranchType = beq & io_IsEq; // @[CU.scala 114:16]
  assign io_IsJType = j | jal; // @[CU.scala 120:14]
  assign io_IsJr = RType & func == 6'h8; // @[CU.scala 86:25]
  assign io_ALUSrc = ori | lui | lw | sw; // @[CU.scala 132:27]
  assign io_WhichToReg = lw ? 2'h1 : _GEN_20; // @[CU.scala 138:23 139:23]
  assign io_RegDst = _T_33 ? 2'h1 : _GEN_20; // @[CU.scala 146:37 147:19]
  assign io_IsSignExt = beq | lw | sw; // @[CU.scala 154:21]
endmodule
module IFU(
  input         clock,
  input         reset,
  input  [31:0] io_NPC,
  output [31:0] io_instr,
  output [31:0] io_PC
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ROM [0:1023]; // @[IFU.scala 12:29]
  wire  ROM_io_instr_MPORT_en; // @[IFU.scala 12:29]
  wire [9:0] ROM_io_instr_MPORT_addr; // @[IFU.scala 12:29]
  wire [31:0] ROM_io_instr_MPORT_data; // @[IFU.scala 12:29]
  reg [31:0] r_PC; // @[IFU.scala 14:19]
  assign ROM_io_instr_MPORT_en = 1'h1;
  assign ROM_io_instr_MPORT_addr = io_PC[11:2];
  assign ROM_io_instr_MPORT_data = ROM[ROM_io_instr_MPORT_addr]; // @[IFU.scala 12:29]
  assign io_instr = ROM_io_instr_MPORT_data; // @[IFU.scala 24:14]
  assign io_PC = r_PC; // @[IFU.scala 23:11]
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 16:25]
      r_PC <= 32'h3000; // @[IFU.scala 19:14]
    end else begin
      r_PC <= io_NPC; // @[IFU.scala 21:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (reset & ~reset) begin
          $fwrite(32'h80000002,"load successfully!"); // @[IFU.scala 18:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
  integer initvar;
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_PC = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
  $readmemh("code.txt", ROM);
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NPC(
  input  [31:0] io_PC,
  input         io_IsBranchType,
  input         io_IsJType,
  input  [31:0] io_instr,
  input         io_IsJr,
  input  [31:0] io_JrAddr,
  input  [31:0] io_imm32,
  output [31:0] io_NPC
);
  wire [31:0] _io_NPC_T_1 = io_PC + 32'h4; // @[NPC.scala 18:25]
  wire [33:0] _GEN_3 = {io_imm32, 2'h0}; // @[NPC.scala 18:43]
  wire [34:0] _io_NPC_T_2 = {{1'd0}, _GEN_3}; // @[NPC.scala 18:43]
  wire [34:0] _GEN_4 = {{3'd0}, _io_NPC_T_1}; // @[NPC.scala 18:31]
  wire [34:0] _io_NPC_T_4 = _GEN_4 + _io_NPC_T_2; // @[NPC.scala 18:31]
  wire [31:0] _io_NPC_T_7 = {io_PC[31:28],io_instr[25:0],2'h0}; // @[Cat.scala 31:58]
  wire [31:0] _GEN_0 = io_IsJr ? io_JrAddr : _io_NPC_T_1; // @[NPC.scala 21:35 22:16 24:16]
  wire [31:0] _GEN_1 = io_IsJType ? _io_NPC_T_7 : _GEN_0; // @[NPC.scala 19:38 20:16]
  wire [34:0] _GEN_2 = io_IsBranchType ? _io_NPC_T_4 : {{3'd0}, _GEN_1}; // @[NPC.scala 17:35 18:16]
  assign io_NPC = _GEN_2[31:0];
endmodule
module GRF(
  input         clock,
  input         reset,
  input  [4:0]  io_A1,
  input  [4:0]  io_A2,
  input  [4:0]  io_A3,
  input         io_WE,
  input  [31:0] io_WD,
  input  [31:0] io_PC,
  output [31:0] io_O1,
  output [31:0] io_O2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_0; // @[GRF.scala 17:29]
  reg [31:0] reg_1; // @[GRF.scala 17:29]
  reg [31:0] reg_2; // @[GRF.scala 17:29]
  reg [31:0] reg_3; // @[GRF.scala 17:29]
  reg [31:0] reg_4; // @[GRF.scala 17:29]
  reg [31:0] reg_5; // @[GRF.scala 17:29]
  reg [31:0] reg_6; // @[GRF.scala 17:29]
  reg [31:0] reg_7; // @[GRF.scala 17:29]
  reg [31:0] reg_8; // @[GRF.scala 17:29]
  reg [31:0] reg_9; // @[GRF.scala 17:29]
  reg [31:0] reg_10; // @[GRF.scala 17:29]
  reg [31:0] reg_11; // @[GRF.scala 17:29]
  reg [31:0] reg_12; // @[GRF.scala 17:29]
  reg [31:0] reg_13; // @[GRF.scala 17:29]
  reg [31:0] reg_14; // @[GRF.scala 17:29]
  reg [31:0] reg_15; // @[GRF.scala 17:29]
  reg [31:0] reg_16; // @[GRF.scala 17:29]
  reg [31:0] reg_17; // @[GRF.scala 17:29]
  reg [31:0] reg_18; // @[GRF.scala 17:29]
  reg [31:0] reg_19; // @[GRF.scala 17:29]
  reg [31:0] reg_20; // @[GRF.scala 17:29]
  reg [31:0] reg_21; // @[GRF.scala 17:29]
  reg [31:0] reg_22; // @[GRF.scala 17:29]
  reg [31:0] reg_23; // @[GRF.scala 17:29]
  reg [31:0] reg_24; // @[GRF.scala 17:29]
  reg [31:0] reg_25; // @[GRF.scala 17:29]
  reg [31:0] reg_26; // @[GRF.scala 17:29]
  reg [31:0] reg_27; // @[GRF.scala 17:29]
  reg [31:0] reg_28; // @[GRF.scala 17:29]
  reg [31:0] reg_29; // @[GRF.scala 17:29]
  reg [31:0] reg_30; // @[GRF.scala 17:29]
  reg [31:0] reg_31; // @[GRF.scala 17:29]
  wire  _T_3 = io_A3 != 5'h0 & io_WE; // @[GRF.scala 22:31]
  wire [31:0] _GEN_97 = 5'h1 == io_A1 ? reg_1 : reg_0; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_98 = 5'h2 == io_A1 ? reg_2 : _GEN_97; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_99 = 5'h3 == io_A1 ? reg_3 : _GEN_98; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_100 = 5'h4 == io_A1 ? reg_4 : _GEN_99; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_101 = 5'h5 == io_A1 ? reg_5 : _GEN_100; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_102 = 5'h6 == io_A1 ? reg_6 : _GEN_101; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_103 = 5'h7 == io_A1 ? reg_7 : _GEN_102; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_104 = 5'h8 == io_A1 ? reg_8 : _GEN_103; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_105 = 5'h9 == io_A1 ? reg_9 : _GEN_104; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_106 = 5'ha == io_A1 ? reg_10 : _GEN_105; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_107 = 5'hb == io_A1 ? reg_11 : _GEN_106; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_108 = 5'hc == io_A1 ? reg_12 : _GEN_107; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_109 = 5'hd == io_A1 ? reg_13 : _GEN_108; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_110 = 5'he == io_A1 ? reg_14 : _GEN_109; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_111 = 5'hf == io_A1 ? reg_15 : _GEN_110; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_112 = 5'h10 == io_A1 ? reg_16 : _GEN_111; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_113 = 5'h11 == io_A1 ? reg_17 : _GEN_112; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_114 = 5'h12 == io_A1 ? reg_18 : _GEN_113; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_115 = 5'h13 == io_A1 ? reg_19 : _GEN_114; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_116 = 5'h14 == io_A1 ? reg_20 : _GEN_115; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_117 = 5'h15 == io_A1 ? reg_21 : _GEN_116; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_118 = 5'h16 == io_A1 ? reg_22 : _GEN_117; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_119 = 5'h17 == io_A1 ? reg_23 : _GEN_118; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_120 = 5'h18 == io_A1 ? reg_24 : _GEN_119; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_121 = 5'h19 == io_A1 ? reg_25 : _GEN_120; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_122 = 5'h1a == io_A1 ? reg_26 : _GEN_121; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_123 = 5'h1b == io_A1 ? reg_27 : _GEN_122; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_124 = 5'h1c == io_A1 ? reg_28 : _GEN_123; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_125 = 5'h1d == io_A1 ? reg_29 : _GEN_124; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_126 = 5'h1e == io_A1 ? reg_30 : _GEN_125; // @[GRF.scala 27:{11,11}]
  wire [31:0] _GEN_129 = 5'h1 == io_A2 ? reg_1 : reg_0; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_130 = 5'h2 == io_A2 ? reg_2 : _GEN_129; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_131 = 5'h3 == io_A2 ? reg_3 : _GEN_130; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_132 = 5'h4 == io_A2 ? reg_4 : _GEN_131; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_133 = 5'h5 == io_A2 ? reg_5 : _GEN_132; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_134 = 5'h6 == io_A2 ? reg_6 : _GEN_133; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_135 = 5'h7 == io_A2 ? reg_7 : _GEN_134; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_136 = 5'h8 == io_A2 ? reg_8 : _GEN_135; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_137 = 5'h9 == io_A2 ? reg_9 : _GEN_136; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_138 = 5'ha == io_A2 ? reg_10 : _GEN_137; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_139 = 5'hb == io_A2 ? reg_11 : _GEN_138; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_140 = 5'hc == io_A2 ? reg_12 : _GEN_139; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_141 = 5'hd == io_A2 ? reg_13 : _GEN_140; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_142 = 5'he == io_A2 ? reg_14 : _GEN_141; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_143 = 5'hf == io_A2 ? reg_15 : _GEN_142; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_144 = 5'h10 == io_A2 ? reg_16 : _GEN_143; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_145 = 5'h11 == io_A2 ? reg_17 : _GEN_144; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_146 = 5'h12 == io_A2 ? reg_18 : _GEN_145; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_147 = 5'h13 == io_A2 ? reg_19 : _GEN_146; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_148 = 5'h14 == io_A2 ? reg_20 : _GEN_147; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_149 = 5'h15 == io_A2 ? reg_21 : _GEN_148; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_150 = 5'h16 == io_A2 ? reg_22 : _GEN_149; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_151 = 5'h17 == io_A2 ? reg_23 : _GEN_150; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_152 = 5'h18 == io_A2 ? reg_24 : _GEN_151; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_153 = 5'h19 == io_A2 ? reg_25 : _GEN_152; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_154 = 5'h1a == io_A2 ? reg_26 : _GEN_153; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_155 = 5'h1b == io_A2 ? reg_27 : _GEN_154; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_156 = 5'h1c == io_A2 ? reg_28 : _GEN_155; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_157 = 5'h1d == io_A2 ? reg_29 : _GEN_156; // @[GRF.scala 28:{11,11}]
  wire [31:0] _GEN_158 = 5'h1e == io_A2 ? reg_30 : _GEN_157; // @[GRF.scala 28:{11,11}]
  assign io_O1 = 5'h1f == io_A1 ? reg_31 : _GEN_126; // @[GRF.scala 27:{11,11}]
  assign io_O2 = 5'h1f == io_A2 ? reg_31 : _GEN_158; // @[GRF.scala 28:{11,11}]
  always @(posedge clock) begin
    if (reset) begin // @[GRF.scala 18:25]
      reg_0 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h0 == io_A3) begin // @[GRF.scala 23:20]
        reg_0 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_1 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h1 == io_A3) begin // @[GRF.scala 23:20]
        reg_1 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_2 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h2 == io_A3) begin // @[GRF.scala 23:20]
        reg_2 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_3 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h3 == io_A3) begin // @[GRF.scala 23:20]
        reg_3 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_4 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h4 == io_A3) begin // @[GRF.scala 23:20]
        reg_4 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_5 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h5 == io_A3) begin // @[GRF.scala 23:20]
        reg_5 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_6 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h6 == io_A3) begin // @[GRF.scala 23:20]
        reg_6 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_7 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h7 == io_A3) begin // @[GRF.scala 23:20]
        reg_7 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_8 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h8 == io_A3) begin // @[GRF.scala 23:20]
        reg_8 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_9 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h9 == io_A3) begin // @[GRF.scala 23:20]
        reg_9 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_10 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'ha == io_A3) begin // @[GRF.scala 23:20]
        reg_10 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_11 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'hb == io_A3) begin // @[GRF.scala 23:20]
        reg_11 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_12 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'hc == io_A3) begin // @[GRF.scala 23:20]
        reg_12 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_13 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'hd == io_A3) begin // @[GRF.scala 23:20]
        reg_13 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_14 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'he == io_A3) begin // @[GRF.scala 23:20]
        reg_14 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_15 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'hf == io_A3) begin // @[GRF.scala 23:20]
        reg_15 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_16 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h10 == io_A3) begin // @[GRF.scala 23:20]
        reg_16 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_17 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h11 == io_A3) begin // @[GRF.scala 23:20]
        reg_17 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_18 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h12 == io_A3) begin // @[GRF.scala 23:20]
        reg_18 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_19 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h13 == io_A3) begin // @[GRF.scala 23:20]
        reg_19 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_20 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h14 == io_A3) begin // @[GRF.scala 23:20]
        reg_20 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_21 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h15 == io_A3) begin // @[GRF.scala 23:20]
        reg_21 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_22 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h16 == io_A3) begin // @[GRF.scala 23:20]
        reg_22 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_23 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h17 == io_A3) begin // @[GRF.scala 23:20]
        reg_23 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_24 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h18 == io_A3) begin // @[GRF.scala 23:20]
        reg_24 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_25 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h19 == io_A3) begin // @[GRF.scala 23:20]
        reg_25 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_26 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h1a == io_A3) begin // @[GRF.scala 23:20]
        reg_26 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_27 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h1b == io_A3) begin // @[GRF.scala 23:20]
        reg_27 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_28 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h1c == io_A3) begin // @[GRF.scala 23:20]
        reg_28 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_29 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h1d == io_A3) begin // @[GRF.scala 23:20]
        reg_29 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_30 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h1e == io_A3) begin // @[GRF.scala 23:20]
        reg_30 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    if (reset) begin // @[GRF.scala 18:25]
      reg_31 <= 32'h0; // @[GRF.scala 20:20]
    end else if (io_A3 != 5'h0 & io_WE) begin // @[GRF.scala 22:49]
      if (5'h1f == io_A3) begin // @[GRF.scala 23:20]
        reg_31 <= io_WD; // @[GRF.scala 23:20]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & _T_3 & ~reset) begin
          $fwrite(32'h80000002,"@0x%x: %d <= 0x%x\n",io_PC,io_A3,io_WD); // @[GRF.scala 24:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  reg_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input  [31:0] io_A1,
  input  [31:0] io_A2,
  input  [3:0]  io_ALUOp,
  output [31:0] io_O,
  output        io_IsEq
);
  wire [31:0] _io_O_T_1 = io_A1 + io_A2; // @[ALU.scala 18:27]
  wire [31:0] _io_O_T_3 = io_A1 - io_A2; // @[ALU.scala 21:27]
  wire [31:0] _io_O_T_4 = io_A1 & io_A2; // @[ALU.scala 24:27]
  wire [31:0] _io_O_T_5 = io_A1 | io_A2; // @[ALU.scala 27:27]
  wire [47:0] _io_O_T_6 = {io_A2, 16'h0}; // @[ALU.scala 30:27]
  wire [47:0] _GEN_0 = 4'h4 == io_ALUOp ? _io_O_T_6 : 48'h0; // @[ALU.scala 15:10 16:23 30:18]
  wire [47:0] _GEN_1 = 4'h3 == io_ALUOp ? {{16'd0}, _io_O_T_5} : _GEN_0; // @[ALU.scala 16:23 27:18]
  wire [47:0] _GEN_2 = 4'h2 == io_ALUOp ? {{16'd0}, _io_O_T_4} : _GEN_1; // @[ALU.scala 16:23 24:18]
  wire [47:0] _GEN_3 = 4'h1 == io_ALUOp ? {{16'd0}, _io_O_T_3} : _GEN_2; // @[ALU.scala 16:23 21:18]
  wire [47:0] _GEN_4 = 4'h0 == io_ALUOp ? {{16'd0}, _io_O_T_1} : _GEN_3; // @[ALU.scala 16:23 18:18]
  assign io_O = _GEN_4[31:0];
  assign io_IsEq = io_A1 == io_A2; // @[ALU.scala 34:17]
endmodule
module DM(
  input         clock,
  input         reset,
  input  [31:0] io_Addr,
  input  [31:0] io_WD,
  input         io_WE,
  input  [31:0] io_PC,
  output [31:0] io_RD
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [31:0] RAM [0:1023]; // @[DM.scala 12:29]
  wire  RAM_io_RD_MPORT_en; // @[DM.scala 12:29]
  wire [9:0] RAM_io_RD_MPORT_addr; // @[DM.scala 12:29]
  wire [31:0] RAM_io_RD_MPORT_data; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_2_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_2_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_2_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_2_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_3_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_3_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_3_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_3_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_4_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_4_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_4_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_4_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_5_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_5_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_5_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_5_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_6_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_6_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_6_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_6_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_7_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_7_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_7_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_7_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_8_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_8_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_8_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_8_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_9_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_9_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_9_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_9_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_10_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_10_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_10_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_10_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_11_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_11_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_11_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_11_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_12_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_12_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_12_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_12_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_13_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_13_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_13_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_13_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_14_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_14_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_14_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_14_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_15_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_15_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_15_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_15_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_16_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_16_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_16_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_16_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_17_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_17_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_17_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_17_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_18_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_18_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_18_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_18_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_19_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_19_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_19_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_19_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_20_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_20_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_20_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_20_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_21_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_21_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_21_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_21_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_22_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_22_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_22_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_22_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_23_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_23_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_23_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_23_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_24_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_24_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_24_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_24_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_25_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_25_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_25_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_25_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_26_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_26_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_26_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_26_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_27_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_27_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_27_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_27_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_28_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_28_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_28_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_28_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_29_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_29_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_29_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_29_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_30_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_30_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_30_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_30_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_31_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_31_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_31_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_31_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_32_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_32_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_32_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_32_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_33_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_33_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_33_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_33_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_34_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_34_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_34_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_34_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_35_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_35_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_35_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_35_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_36_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_36_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_36_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_36_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_37_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_37_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_37_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_37_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_38_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_38_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_38_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_38_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_39_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_39_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_39_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_39_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_40_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_40_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_40_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_40_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_41_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_41_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_41_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_41_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_42_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_42_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_42_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_42_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_43_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_43_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_43_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_43_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_44_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_44_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_44_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_44_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_45_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_45_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_45_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_45_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_46_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_46_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_46_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_46_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_47_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_47_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_47_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_47_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_48_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_48_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_48_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_48_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_49_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_49_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_49_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_49_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_50_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_50_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_50_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_50_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_51_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_51_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_51_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_51_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_52_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_52_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_52_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_52_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_53_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_53_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_53_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_53_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_54_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_54_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_54_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_54_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_55_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_55_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_55_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_55_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_56_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_56_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_56_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_56_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_57_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_57_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_57_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_57_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_58_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_58_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_58_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_58_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_59_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_59_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_59_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_59_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_60_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_60_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_60_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_60_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_61_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_61_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_61_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_61_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_62_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_62_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_62_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_62_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_63_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_63_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_63_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_63_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_64_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_64_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_64_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_64_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_65_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_65_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_65_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_65_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_66_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_66_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_66_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_66_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_67_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_67_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_67_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_67_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_68_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_68_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_68_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_68_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_69_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_69_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_69_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_69_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_70_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_70_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_70_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_70_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_71_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_71_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_71_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_71_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_72_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_72_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_72_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_72_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_73_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_73_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_73_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_73_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_74_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_74_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_74_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_74_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_75_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_75_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_75_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_75_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_76_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_76_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_76_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_76_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_77_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_77_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_77_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_77_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_78_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_78_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_78_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_78_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_79_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_79_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_79_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_79_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_80_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_80_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_80_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_80_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_81_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_81_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_81_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_81_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_82_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_82_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_82_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_82_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_83_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_83_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_83_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_83_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_84_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_84_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_84_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_84_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_85_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_85_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_85_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_85_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_86_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_86_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_86_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_86_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_87_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_87_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_87_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_87_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_88_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_88_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_88_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_88_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_89_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_89_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_89_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_89_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_90_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_90_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_90_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_90_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_91_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_91_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_91_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_91_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_92_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_92_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_92_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_92_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_93_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_93_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_93_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_93_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_94_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_94_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_94_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_94_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_95_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_95_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_95_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_95_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_96_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_96_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_96_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_96_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_97_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_97_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_97_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_97_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_98_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_98_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_98_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_98_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_99_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_99_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_99_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_99_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_100_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_100_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_100_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_100_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_101_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_101_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_101_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_101_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_102_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_102_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_102_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_102_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_103_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_103_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_103_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_103_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_104_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_104_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_104_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_104_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_105_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_105_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_105_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_105_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_106_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_106_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_106_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_106_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_107_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_107_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_107_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_107_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_108_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_108_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_108_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_108_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_109_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_109_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_109_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_109_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_110_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_110_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_110_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_110_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_111_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_111_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_111_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_111_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_112_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_112_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_112_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_112_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_113_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_113_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_113_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_113_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_114_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_114_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_114_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_114_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_115_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_115_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_115_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_115_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_116_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_116_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_116_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_116_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_117_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_117_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_117_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_117_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_118_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_118_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_118_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_118_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_119_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_119_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_119_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_119_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_120_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_120_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_120_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_120_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_121_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_121_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_121_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_121_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_122_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_122_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_122_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_122_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_123_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_123_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_123_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_123_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_124_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_124_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_124_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_124_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_125_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_125_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_125_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_125_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_126_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_126_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_126_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_126_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_127_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_127_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_127_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_127_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_128_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_128_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_128_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_128_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_129_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_129_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_129_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_129_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_130_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_130_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_130_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_130_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_131_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_131_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_131_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_131_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_132_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_132_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_132_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_132_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_133_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_133_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_133_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_133_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_134_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_134_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_134_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_134_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_135_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_135_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_135_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_135_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_136_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_136_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_136_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_136_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_137_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_137_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_137_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_137_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_138_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_138_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_138_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_138_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_139_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_139_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_139_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_139_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_140_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_140_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_140_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_140_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_141_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_141_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_141_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_141_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_142_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_142_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_142_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_142_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_143_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_143_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_143_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_143_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_144_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_144_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_144_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_144_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_145_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_145_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_145_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_145_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_146_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_146_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_146_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_146_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_147_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_147_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_147_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_147_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_148_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_148_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_148_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_148_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_149_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_149_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_149_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_149_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_150_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_150_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_150_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_150_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_151_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_151_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_151_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_151_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_152_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_152_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_152_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_152_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_153_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_153_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_153_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_153_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_154_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_154_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_154_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_154_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_155_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_155_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_155_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_155_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_156_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_156_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_156_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_156_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_157_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_157_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_157_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_157_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_158_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_158_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_158_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_158_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_159_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_159_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_159_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_159_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_160_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_160_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_160_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_160_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_161_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_161_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_161_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_161_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_162_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_162_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_162_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_162_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_163_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_163_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_163_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_163_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_164_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_164_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_164_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_164_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_165_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_165_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_165_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_165_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_166_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_166_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_166_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_166_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_167_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_167_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_167_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_167_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_168_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_168_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_168_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_168_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_169_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_169_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_169_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_169_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_170_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_170_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_170_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_170_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_171_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_171_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_171_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_171_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_172_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_172_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_172_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_172_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_173_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_173_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_173_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_173_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_174_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_174_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_174_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_174_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_175_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_175_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_175_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_175_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_176_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_176_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_176_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_176_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_177_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_177_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_177_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_177_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_178_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_178_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_178_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_178_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_179_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_179_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_179_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_179_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_180_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_180_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_180_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_180_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_181_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_181_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_181_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_181_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_182_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_182_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_182_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_182_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_183_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_183_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_183_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_183_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_184_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_184_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_184_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_184_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_185_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_185_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_185_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_185_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_186_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_186_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_186_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_186_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_187_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_187_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_187_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_187_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_188_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_188_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_188_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_188_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_189_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_189_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_189_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_189_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_190_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_190_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_190_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_190_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_191_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_191_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_191_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_191_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_192_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_192_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_192_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_192_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_193_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_193_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_193_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_193_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_194_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_194_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_194_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_194_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_195_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_195_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_195_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_195_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_196_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_196_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_196_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_196_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_197_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_197_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_197_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_197_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_198_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_198_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_198_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_198_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_199_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_199_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_199_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_199_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_200_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_200_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_200_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_200_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_201_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_201_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_201_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_201_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_202_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_202_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_202_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_202_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_203_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_203_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_203_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_203_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_204_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_204_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_204_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_204_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_205_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_205_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_205_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_205_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_206_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_206_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_206_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_206_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_207_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_207_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_207_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_207_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_208_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_208_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_208_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_208_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_209_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_209_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_209_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_209_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_210_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_210_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_210_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_210_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_211_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_211_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_211_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_211_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_212_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_212_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_212_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_212_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_213_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_213_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_213_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_213_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_214_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_214_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_214_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_214_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_215_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_215_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_215_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_215_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_216_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_216_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_216_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_216_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_217_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_217_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_217_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_217_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_218_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_218_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_218_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_218_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_219_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_219_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_219_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_219_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_220_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_220_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_220_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_220_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_221_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_221_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_221_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_221_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_222_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_222_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_222_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_222_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_223_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_223_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_223_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_223_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_224_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_224_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_224_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_224_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_225_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_225_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_225_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_225_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_226_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_226_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_226_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_226_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_227_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_227_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_227_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_227_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_228_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_228_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_228_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_228_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_229_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_229_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_229_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_229_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_230_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_230_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_230_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_230_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_231_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_231_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_231_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_231_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_232_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_232_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_232_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_232_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_233_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_233_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_233_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_233_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_234_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_234_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_234_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_234_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_235_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_235_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_235_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_235_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_236_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_236_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_236_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_236_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_237_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_237_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_237_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_237_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_238_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_238_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_238_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_238_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_239_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_239_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_239_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_239_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_240_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_240_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_240_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_240_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_241_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_241_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_241_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_241_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_242_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_242_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_242_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_242_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_243_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_243_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_243_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_243_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_244_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_244_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_244_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_244_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_245_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_245_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_245_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_245_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_246_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_246_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_246_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_246_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_247_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_247_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_247_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_247_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_248_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_248_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_248_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_248_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_249_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_249_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_249_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_249_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_250_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_250_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_250_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_250_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_251_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_251_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_251_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_251_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_252_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_252_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_252_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_252_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_253_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_253_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_253_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_253_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_254_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_254_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_254_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_254_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_255_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_255_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_255_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_255_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_256_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_256_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_256_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_256_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_257_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_257_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_257_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_257_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_258_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_258_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_258_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_258_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_259_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_259_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_259_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_259_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_260_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_260_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_260_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_260_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_261_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_261_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_261_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_261_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_262_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_262_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_262_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_262_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_263_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_263_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_263_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_263_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_264_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_264_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_264_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_264_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_265_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_265_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_265_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_265_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_266_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_266_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_266_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_266_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_267_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_267_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_267_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_267_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_268_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_268_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_268_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_268_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_269_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_269_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_269_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_269_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_270_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_270_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_270_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_270_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_271_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_271_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_271_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_271_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_272_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_272_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_272_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_272_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_273_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_273_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_273_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_273_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_274_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_274_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_274_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_274_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_275_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_275_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_275_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_275_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_276_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_276_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_276_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_276_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_277_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_277_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_277_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_277_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_278_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_278_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_278_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_278_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_279_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_279_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_279_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_279_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_280_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_280_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_280_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_280_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_281_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_281_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_281_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_281_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_282_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_282_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_282_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_282_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_283_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_283_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_283_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_283_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_284_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_284_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_284_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_284_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_285_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_285_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_285_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_285_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_286_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_286_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_286_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_286_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_287_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_287_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_287_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_287_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_288_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_288_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_288_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_288_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_289_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_289_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_289_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_289_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_290_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_290_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_290_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_290_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_291_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_291_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_291_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_291_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_292_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_292_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_292_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_292_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_293_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_293_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_293_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_293_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_294_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_294_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_294_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_294_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_295_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_295_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_295_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_295_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_296_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_296_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_296_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_296_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_297_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_297_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_297_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_297_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_298_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_298_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_298_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_298_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_299_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_299_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_299_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_299_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_300_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_300_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_300_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_300_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_301_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_301_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_301_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_301_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_302_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_302_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_302_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_302_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_303_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_303_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_303_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_303_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_304_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_304_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_304_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_304_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_305_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_305_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_305_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_305_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_306_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_306_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_306_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_306_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_307_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_307_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_307_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_307_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_308_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_308_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_308_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_308_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_309_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_309_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_309_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_309_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_310_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_310_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_310_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_310_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_311_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_311_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_311_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_311_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_312_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_312_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_312_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_312_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_313_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_313_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_313_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_313_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_314_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_314_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_314_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_314_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_315_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_315_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_315_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_315_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_316_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_316_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_316_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_316_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_317_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_317_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_317_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_317_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_318_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_318_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_318_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_318_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_319_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_319_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_319_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_319_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_320_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_320_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_320_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_320_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_321_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_321_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_321_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_321_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_322_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_322_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_322_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_322_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_323_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_323_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_323_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_323_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_324_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_324_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_324_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_324_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_325_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_325_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_325_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_325_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_326_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_326_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_326_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_326_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_327_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_327_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_327_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_327_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_328_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_328_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_328_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_328_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_329_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_329_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_329_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_329_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_330_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_330_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_330_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_330_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_331_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_331_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_331_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_331_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_332_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_332_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_332_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_332_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_333_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_333_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_333_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_333_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_334_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_334_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_334_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_334_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_335_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_335_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_335_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_335_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_336_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_336_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_336_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_336_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_337_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_337_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_337_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_337_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_338_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_338_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_338_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_338_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_339_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_339_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_339_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_339_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_340_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_340_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_340_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_340_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_341_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_341_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_341_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_341_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_342_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_342_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_342_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_342_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_343_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_343_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_343_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_343_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_344_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_344_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_344_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_344_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_345_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_345_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_345_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_345_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_346_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_346_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_346_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_346_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_347_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_347_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_347_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_347_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_348_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_348_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_348_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_348_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_349_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_349_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_349_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_349_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_350_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_350_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_350_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_350_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_351_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_351_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_351_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_351_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_352_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_352_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_352_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_352_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_353_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_353_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_353_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_353_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_354_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_354_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_354_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_354_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_355_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_355_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_355_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_355_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_356_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_356_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_356_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_356_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_357_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_357_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_357_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_357_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_358_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_358_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_358_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_358_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_359_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_359_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_359_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_359_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_360_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_360_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_360_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_360_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_361_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_361_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_361_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_361_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_362_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_362_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_362_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_362_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_363_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_363_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_363_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_363_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_364_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_364_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_364_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_364_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_365_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_365_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_365_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_365_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_366_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_366_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_366_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_366_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_367_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_367_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_367_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_367_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_368_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_368_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_368_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_368_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_369_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_369_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_369_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_369_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_370_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_370_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_370_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_370_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_371_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_371_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_371_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_371_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_372_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_372_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_372_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_372_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_373_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_373_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_373_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_373_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_374_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_374_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_374_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_374_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_375_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_375_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_375_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_375_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_376_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_376_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_376_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_376_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_377_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_377_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_377_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_377_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_378_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_378_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_378_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_378_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_379_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_379_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_379_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_379_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_380_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_380_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_380_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_380_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_381_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_381_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_381_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_381_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_382_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_382_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_382_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_382_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_383_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_383_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_383_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_383_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_384_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_384_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_384_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_384_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_385_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_385_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_385_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_385_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_386_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_386_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_386_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_386_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_387_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_387_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_387_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_387_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_388_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_388_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_388_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_388_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_389_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_389_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_389_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_389_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_390_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_390_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_390_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_390_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_391_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_391_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_391_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_391_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_392_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_392_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_392_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_392_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_393_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_393_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_393_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_393_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_394_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_394_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_394_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_394_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_395_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_395_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_395_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_395_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_396_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_396_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_396_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_396_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_397_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_397_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_397_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_397_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_398_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_398_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_398_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_398_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_399_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_399_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_399_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_399_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_400_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_400_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_400_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_400_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_401_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_401_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_401_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_401_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_402_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_402_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_402_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_402_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_403_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_403_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_403_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_403_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_404_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_404_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_404_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_404_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_405_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_405_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_405_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_405_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_406_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_406_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_406_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_406_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_407_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_407_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_407_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_407_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_408_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_408_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_408_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_408_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_409_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_409_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_409_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_409_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_410_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_410_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_410_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_410_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_411_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_411_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_411_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_411_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_412_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_412_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_412_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_412_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_413_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_413_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_413_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_413_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_414_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_414_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_414_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_414_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_415_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_415_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_415_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_415_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_416_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_416_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_416_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_416_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_417_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_417_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_417_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_417_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_418_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_418_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_418_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_418_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_419_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_419_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_419_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_419_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_420_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_420_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_420_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_420_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_421_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_421_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_421_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_421_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_422_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_422_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_422_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_422_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_423_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_423_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_423_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_423_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_424_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_424_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_424_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_424_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_425_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_425_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_425_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_425_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_426_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_426_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_426_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_426_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_427_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_427_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_427_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_427_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_428_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_428_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_428_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_428_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_429_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_429_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_429_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_429_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_430_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_430_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_430_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_430_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_431_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_431_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_431_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_431_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_432_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_432_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_432_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_432_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_433_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_433_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_433_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_433_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_434_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_434_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_434_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_434_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_435_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_435_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_435_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_435_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_436_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_436_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_436_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_436_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_437_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_437_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_437_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_437_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_438_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_438_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_438_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_438_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_439_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_439_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_439_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_439_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_440_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_440_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_440_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_440_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_441_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_441_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_441_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_441_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_442_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_442_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_442_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_442_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_443_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_443_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_443_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_443_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_444_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_444_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_444_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_444_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_445_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_445_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_445_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_445_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_446_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_446_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_446_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_446_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_447_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_447_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_447_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_447_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_448_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_448_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_448_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_448_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_449_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_449_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_449_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_449_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_450_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_450_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_450_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_450_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_451_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_451_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_451_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_451_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_452_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_452_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_452_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_452_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_453_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_453_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_453_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_453_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_454_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_454_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_454_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_454_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_455_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_455_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_455_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_455_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_456_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_456_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_456_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_456_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_457_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_457_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_457_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_457_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_458_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_458_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_458_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_458_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_459_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_459_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_459_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_459_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_460_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_460_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_460_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_460_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_461_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_461_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_461_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_461_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_462_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_462_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_462_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_462_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_463_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_463_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_463_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_463_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_464_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_464_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_464_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_464_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_465_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_465_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_465_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_465_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_466_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_466_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_466_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_466_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_467_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_467_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_467_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_467_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_468_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_468_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_468_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_468_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_469_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_469_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_469_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_469_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_470_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_470_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_470_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_470_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_471_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_471_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_471_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_471_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_472_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_472_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_472_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_472_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_473_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_473_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_473_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_473_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_474_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_474_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_474_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_474_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_475_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_475_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_475_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_475_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_476_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_476_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_476_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_476_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_477_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_477_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_477_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_477_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_478_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_478_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_478_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_478_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_479_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_479_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_479_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_479_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_480_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_480_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_480_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_480_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_481_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_481_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_481_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_481_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_482_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_482_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_482_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_482_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_483_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_483_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_483_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_483_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_484_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_484_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_484_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_484_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_485_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_485_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_485_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_485_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_486_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_486_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_486_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_486_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_487_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_487_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_487_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_487_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_488_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_488_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_488_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_488_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_489_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_489_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_489_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_489_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_490_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_490_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_490_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_490_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_491_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_491_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_491_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_491_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_492_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_492_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_492_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_492_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_493_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_493_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_493_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_493_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_494_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_494_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_494_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_494_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_495_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_495_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_495_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_495_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_496_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_496_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_496_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_496_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_497_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_497_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_497_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_497_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_498_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_498_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_498_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_498_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_499_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_499_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_499_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_499_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_500_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_500_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_500_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_500_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_501_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_501_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_501_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_501_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_502_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_502_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_502_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_502_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_503_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_503_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_503_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_503_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_504_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_504_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_504_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_504_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_505_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_505_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_505_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_505_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_506_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_506_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_506_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_506_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_507_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_507_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_507_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_507_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_508_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_508_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_508_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_508_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_509_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_509_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_509_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_509_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_510_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_510_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_510_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_510_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_511_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_511_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_511_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_511_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_512_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_512_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_512_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_512_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_513_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_513_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_513_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_513_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_514_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_514_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_514_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_514_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_515_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_515_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_515_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_515_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_516_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_516_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_516_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_516_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_517_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_517_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_517_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_517_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_518_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_518_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_518_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_518_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_519_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_519_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_519_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_519_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_520_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_520_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_520_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_520_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_521_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_521_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_521_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_521_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_522_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_522_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_522_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_522_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_523_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_523_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_523_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_523_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_524_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_524_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_524_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_524_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_525_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_525_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_525_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_525_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_526_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_526_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_526_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_526_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_527_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_527_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_527_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_527_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_528_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_528_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_528_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_528_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_529_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_529_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_529_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_529_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_530_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_530_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_530_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_530_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_531_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_531_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_531_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_531_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_532_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_532_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_532_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_532_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_533_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_533_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_533_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_533_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_534_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_534_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_534_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_534_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_535_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_535_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_535_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_535_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_536_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_536_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_536_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_536_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_537_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_537_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_537_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_537_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_538_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_538_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_538_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_538_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_539_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_539_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_539_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_539_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_540_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_540_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_540_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_540_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_541_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_541_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_541_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_541_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_542_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_542_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_542_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_542_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_543_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_543_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_543_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_543_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_544_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_544_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_544_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_544_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_545_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_545_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_545_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_545_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_546_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_546_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_546_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_546_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_547_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_547_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_547_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_547_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_548_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_548_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_548_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_548_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_549_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_549_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_549_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_549_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_550_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_550_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_550_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_550_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_551_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_551_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_551_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_551_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_552_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_552_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_552_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_552_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_553_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_553_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_553_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_553_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_554_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_554_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_554_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_554_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_555_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_555_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_555_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_555_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_556_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_556_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_556_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_556_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_557_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_557_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_557_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_557_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_558_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_558_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_558_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_558_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_559_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_559_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_559_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_559_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_560_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_560_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_560_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_560_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_561_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_561_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_561_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_561_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_562_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_562_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_562_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_562_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_563_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_563_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_563_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_563_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_564_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_564_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_564_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_564_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_565_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_565_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_565_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_565_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_566_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_566_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_566_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_566_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_567_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_567_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_567_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_567_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_568_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_568_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_568_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_568_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_569_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_569_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_569_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_569_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_570_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_570_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_570_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_570_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_571_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_571_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_571_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_571_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_572_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_572_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_572_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_572_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_573_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_573_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_573_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_573_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_574_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_574_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_574_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_574_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_575_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_575_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_575_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_575_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_576_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_576_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_576_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_576_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_577_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_577_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_577_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_577_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_578_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_578_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_578_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_578_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_579_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_579_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_579_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_579_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_580_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_580_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_580_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_580_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_581_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_581_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_581_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_581_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_582_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_582_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_582_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_582_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_583_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_583_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_583_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_583_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_584_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_584_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_584_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_584_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_585_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_585_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_585_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_585_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_586_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_586_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_586_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_586_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_587_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_587_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_587_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_587_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_588_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_588_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_588_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_588_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_589_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_589_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_589_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_589_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_590_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_590_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_590_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_590_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_591_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_591_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_591_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_591_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_592_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_592_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_592_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_592_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_593_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_593_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_593_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_593_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_594_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_594_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_594_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_594_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_595_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_595_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_595_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_595_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_596_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_596_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_596_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_596_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_597_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_597_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_597_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_597_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_598_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_598_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_598_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_598_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_599_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_599_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_599_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_599_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_600_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_600_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_600_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_600_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_601_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_601_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_601_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_601_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_602_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_602_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_602_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_602_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_603_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_603_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_603_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_603_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_604_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_604_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_604_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_604_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_605_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_605_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_605_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_605_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_606_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_606_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_606_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_606_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_607_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_607_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_607_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_607_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_608_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_608_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_608_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_608_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_609_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_609_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_609_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_609_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_610_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_610_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_610_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_610_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_611_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_611_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_611_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_611_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_612_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_612_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_612_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_612_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_613_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_613_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_613_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_613_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_614_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_614_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_614_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_614_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_615_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_615_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_615_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_615_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_616_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_616_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_616_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_616_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_617_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_617_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_617_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_617_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_618_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_618_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_618_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_618_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_619_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_619_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_619_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_619_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_620_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_620_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_620_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_620_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_621_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_621_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_621_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_621_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_622_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_622_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_622_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_622_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_623_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_623_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_623_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_623_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_624_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_624_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_624_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_624_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_625_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_625_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_625_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_625_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_626_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_626_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_626_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_626_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_627_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_627_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_627_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_627_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_628_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_628_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_628_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_628_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_629_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_629_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_629_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_629_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_630_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_630_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_630_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_630_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_631_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_631_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_631_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_631_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_632_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_632_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_632_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_632_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_633_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_633_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_633_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_633_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_634_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_634_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_634_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_634_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_635_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_635_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_635_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_635_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_636_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_636_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_636_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_636_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_637_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_637_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_637_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_637_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_638_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_638_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_638_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_638_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_639_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_639_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_639_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_639_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_640_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_640_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_640_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_640_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_641_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_641_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_641_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_641_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_642_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_642_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_642_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_642_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_643_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_643_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_643_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_643_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_644_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_644_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_644_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_644_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_645_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_645_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_645_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_645_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_646_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_646_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_646_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_646_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_647_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_647_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_647_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_647_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_648_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_648_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_648_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_648_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_649_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_649_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_649_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_649_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_650_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_650_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_650_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_650_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_651_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_651_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_651_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_651_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_652_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_652_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_652_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_652_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_653_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_653_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_653_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_653_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_654_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_654_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_654_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_654_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_655_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_655_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_655_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_655_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_656_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_656_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_656_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_656_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_657_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_657_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_657_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_657_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_658_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_658_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_658_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_658_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_659_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_659_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_659_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_659_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_660_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_660_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_660_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_660_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_661_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_661_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_661_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_661_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_662_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_662_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_662_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_662_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_663_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_663_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_663_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_663_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_664_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_664_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_664_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_664_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_665_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_665_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_665_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_665_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_666_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_666_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_666_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_666_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_667_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_667_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_667_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_667_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_668_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_668_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_668_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_668_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_669_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_669_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_669_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_669_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_670_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_670_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_670_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_670_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_671_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_671_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_671_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_671_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_672_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_672_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_672_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_672_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_673_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_673_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_673_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_673_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_674_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_674_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_674_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_674_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_675_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_675_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_675_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_675_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_676_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_676_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_676_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_676_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_677_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_677_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_677_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_677_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_678_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_678_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_678_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_678_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_679_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_679_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_679_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_679_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_680_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_680_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_680_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_680_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_681_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_681_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_681_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_681_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_682_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_682_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_682_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_682_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_683_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_683_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_683_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_683_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_684_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_684_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_684_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_684_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_685_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_685_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_685_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_685_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_686_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_686_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_686_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_686_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_687_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_687_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_687_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_687_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_688_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_688_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_688_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_688_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_689_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_689_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_689_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_689_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_690_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_690_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_690_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_690_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_691_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_691_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_691_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_691_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_692_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_692_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_692_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_692_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_693_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_693_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_693_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_693_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_694_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_694_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_694_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_694_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_695_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_695_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_695_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_695_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_696_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_696_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_696_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_696_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_697_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_697_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_697_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_697_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_698_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_698_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_698_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_698_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_699_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_699_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_699_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_699_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_700_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_700_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_700_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_700_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_701_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_701_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_701_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_701_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_702_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_702_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_702_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_702_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_703_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_703_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_703_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_703_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_704_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_704_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_704_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_704_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_705_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_705_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_705_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_705_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_706_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_706_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_706_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_706_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_707_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_707_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_707_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_707_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_708_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_708_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_708_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_708_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_709_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_709_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_709_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_709_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_710_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_710_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_710_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_710_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_711_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_711_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_711_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_711_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_712_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_712_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_712_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_712_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_713_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_713_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_713_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_713_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_714_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_714_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_714_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_714_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_715_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_715_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_715_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_715_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_716_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_716_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_716_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_716_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_717_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_717_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_717_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_717_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_718_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_718_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_718_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_718_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_719_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_719_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_719_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_719_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_720_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_720_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_720_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_720_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_721_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_721_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_721_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_721_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_722_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_722_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_722_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_722_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_723_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_723_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_723_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_723_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_724_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_724_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_724_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_724_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_725_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_725_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_725_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_725_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_726_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_726_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_726_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_726_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_727_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_727_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_727_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_727_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_728_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_728_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_728_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_728_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_729_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_729_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_729_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_729_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_730_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_730_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_730_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_730_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_731_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_731_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_731_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_731_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_732_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_732_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_732_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_732_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_733_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_733_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_733_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_733_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_734_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_734_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_734_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_734_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_735_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_735_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_735_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_735_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_736_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_736_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_736_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_736_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_737_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_737_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_737_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_737_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_738_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_738_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_738_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_738_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_739_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_739_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_739_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_739_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_740_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_740_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_740_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_740_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_741_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_741_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_741_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_741_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_742_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_742_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_742_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_742_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_743_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_743_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_743_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_743_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_744_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_744_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_744_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_744_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_745_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_745_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_745_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_745_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_746_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_746_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_746_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_746_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_747_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_747_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_747_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_747_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_748_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_748_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_748_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_748_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_749_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_749_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_749_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_749_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_750_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_750_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_750_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_750_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_751_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_751_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_751_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_751_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_752_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_752_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_752_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_752_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_753_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_753_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_753_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_753_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_754_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_754_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_754_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_754_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_755_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_755_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_755_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_755_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_756_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_756_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_756_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_756_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_757_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_757_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_757_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_757_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_758_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_758_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_758_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_758_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_759_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_759_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_759_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_759_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_760_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_760_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_760_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_760_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_761_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_761_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_761_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_761_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_762_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_762_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_762_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_762_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_763_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_763_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_763_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_763_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_764_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_764_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_764_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_764_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_765_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_765_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_765_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_765_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_766_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_766_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_766_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_766_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_767_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_767_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_767_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_767_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_768_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_768_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_768_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_768_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_769_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_769_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_769_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_769_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_770_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_770_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_770_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_770_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_771_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_771_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_771_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_771_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_772_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_772_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_772_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_772_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_773_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_773_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_773_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_773_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_774_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_774_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_774_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_774_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_775_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_775_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_775_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_775_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_776_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_776_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_776_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_776_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_777_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_777_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_777_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_777_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_778_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_778_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_778_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_778_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_779_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_779_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_779_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_779_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_780_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_780_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_780_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_780_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_781_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_781_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_781_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_781_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_782_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_782_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_782_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_782_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_783_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_783_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_783_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_783_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_784_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_784_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_784_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_784_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_785_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_785_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_785_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_785_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_786_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_786_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_786_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_786_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_787_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_787_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_787_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_787_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_788_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_788_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_788_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_788_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_789_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_789_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_789_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_789_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_790_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_790_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_790_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_790_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_791_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_791_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_791_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_791_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_792_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_792_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_792_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_792_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_793_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_793_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_793_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_793_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_794_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_794_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_794_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_794_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_795_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_795_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_795_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_795_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_796_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_796_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_796_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_796_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_797_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_797_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_797_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_797_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_798_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_798_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_798_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_798_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_799_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_799_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_799_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_799_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_800_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_800_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_800_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_800_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_801_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_801_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_801_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_801_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_802_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_802_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_802_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_802_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_803_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_803_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_803_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_803_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_804_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_804_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_804_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_804_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_805_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_805_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_805_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_805_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_806_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_806_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_806_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_806_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_807_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_807_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_807_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_807_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_808_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_808_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_808_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_808_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_809_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_809_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_809_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_809_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_810_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_810_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_810_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_810_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_811_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_811_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_811_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_811_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_812_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_812_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_812_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_812_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_813_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_813_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_813_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_813_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_814_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_814_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_814_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_814_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_815_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_815_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_815_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_815_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_816_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_816_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_816_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_816_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_817_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_817_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_817_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_817_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_818_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_818_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_818_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_818_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_819_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_819_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_819_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_819_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_820_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_820_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_820_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_820_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_821_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_821_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_821_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_821_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_822_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_822_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_822_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_822_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_823_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_823_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_823_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_823_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_824_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_824_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_824_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_824_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_825_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_825_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_825_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_825_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_826_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_826_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_826_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_826_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_827_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_827_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_827_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_827_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_828_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_828_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_828_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_828_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_829_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_829_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_829_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_829_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_830_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_830_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_830_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_830_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_831_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_831_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_831_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_831_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_832_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_832_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_832_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_832_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_833_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_833_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_833_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_833_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_834_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_834_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_834_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_834_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_835_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_835_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_835_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_835_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_836_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_836_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_836_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_836_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_837_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_837_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_837_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_837_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_838_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_838_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_838_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_838_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_839_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_839_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_839_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_839_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_840_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_840_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_840_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_840_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_841_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_841_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_841_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_841_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_842_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_842_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_842_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_842_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_843_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_843_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_843_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_843_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_844_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_844_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_844_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_844_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_845_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_845_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_845_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_845_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_846_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_846_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_846_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_846_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_847_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_847_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_847_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_847_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_848_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_848_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_848_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_848_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_849_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_849_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_849_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_849_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_850_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_850_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_850_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_850_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_851_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_851_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_851_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_851_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_852_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_852_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_852_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_852_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_853_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_853_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_853_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_853_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_854_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_854_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_854_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_854_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_855_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_855_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_855_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_855_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_856_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_856_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_856_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_856_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_857_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_857_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_857_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_857_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_858_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_858_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_858_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_858_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_859_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_859_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_859_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_859_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_860_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_860_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_860_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_860_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_861_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_861_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_861_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_861_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_862_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_862_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_862_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_862_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_863_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_863_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_863_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_863_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_864_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_864_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_864_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_864_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_865_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_865_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_865_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_865_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_866_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_866_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_866_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_866_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_867_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_867_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_867_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_867_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_868_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_868_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_868_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_868_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_869_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_869_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_869_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_869_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_870_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_870_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_870_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_870_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_871_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_871_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_871_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_871_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_872_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_872_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_872_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_872_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_873_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_873_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_873_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_873_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_874_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_874_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_874_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_874_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_875_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_875_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_875_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_875_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_876_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_876_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_876_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_876_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_877_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_877_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_877_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_877_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_878_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_878_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_878_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_878_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_879_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_879_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_879_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_879_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_880_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_880_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_880_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_880_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_881_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_881_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_881_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_881_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_882_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_882_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_882_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_882_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_883_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_883_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_883_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_883_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_884_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_884_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_884_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_884_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_885_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_885_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_885_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_885_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_886_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_886_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_886_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_886_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_887_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_887_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_887_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_887_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_888_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_888_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_888_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_888_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_889_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_889_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_889_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_889_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_890_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_890_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_890_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_890_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_891_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_891_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_891_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_891_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_892_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_892_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_892_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_892_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_893_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_893_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_893_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_893_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_894_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_894_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_894_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_894_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_895_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_895_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_895_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_895_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_896_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_896_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_896_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_896_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_897_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_897_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_897_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_897_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_898_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_898_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_898_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_898_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_899_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_899_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_899_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_899_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_900_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_900_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_900_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_900_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_901_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_901_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_901_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_901_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_902_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_902_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_902_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_902_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_903_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_903_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_903_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_903_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_904_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_904_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_904_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_904_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_905_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_905_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_905_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_905_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_906_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_906_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_906_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_906_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_907_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_907_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_907_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_907_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_908_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_908_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_908_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_908_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_909_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_909_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_909_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_909_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_910_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_910_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_910_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_910_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_911_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_911_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_911_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_911_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_912_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_912_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_912_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_912_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_913_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_913_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_913_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_913_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_914_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_914_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_914_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_914_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_915_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_915_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_915_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_915_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_916_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_916_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_916_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_916_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_917_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_917_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_917_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_917_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_918_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_918_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_918_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_918_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_919_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_919_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_919_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_919_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_920_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_920_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_920_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_920_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_921_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_921_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_921_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_921_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_922_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_922_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_922_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_922_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_923_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_923_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_923_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_923_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_924_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_924_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_924_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_924_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_925_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_925_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_925_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_925_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_926_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_926_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_926_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_926_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_927_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_927_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_927_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_927_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_928_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_928_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_928_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_928_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_929_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_929_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_929_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_929_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_930_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_930_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_930_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_930_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_931_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_931_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_931_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_931_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_932_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_932_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_932_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_932_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_933_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_933_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_933_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_933_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_934_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_934_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_934_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_934_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_935_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_935_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_935_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_935_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_936_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_936_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_936_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_936_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_937_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_937_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_937_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_937_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_938_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_938_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_938_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_938_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_939_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_939_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_939_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_939_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_940_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_940_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_940_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_940_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_941_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_941_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_941_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_941_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_942_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_942_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_942_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_942_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_943_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_943_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_943_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_943_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_944_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_944_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_944_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_944_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_945_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_945_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_945_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_945_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_946_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_946_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_946_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_946_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_947_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_947_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_947_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_947_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_948_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_948_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_948_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_948_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_949_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_949_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_949_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_949_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_950_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_950_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_950_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_950_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_951_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_951_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_951_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_951_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_952_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_952_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_952_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_952_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_953_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_953_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_953_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_953_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_954_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_954_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_954_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_954_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_955_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_955_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_955_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_955_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_956_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_956_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_956_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_956_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_957_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_957_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_957_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_957_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_958_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_958_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_958_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_958_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_959_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_959_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_959_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_959_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_960_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_960_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_960_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_960_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_961_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_961_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_961_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_961_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_962_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_962_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_962_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_962_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_963_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_963_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_963_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_963_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_964_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_964_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_964_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_964_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_965_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_965_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_965_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_965_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_966_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_966_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_966_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_966_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_967_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_967_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_967_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_967_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_968_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_968_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_968_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_968_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_969_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_969_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_969_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_969_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_970_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_970_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_970_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_970_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_971_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_971_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_971_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_971_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_972_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_972_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_972_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_972_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_973_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_973_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_973_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_973_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_974_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_974_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_974_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_974_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_975_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_975_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_975_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_975_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_976_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_976_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_976_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_976_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_977_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_977_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_977_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_977_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_978_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_978_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_978_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_978_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_979_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_979_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_979_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_979_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_980_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_980_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_980_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_980_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_981_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_981_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_981_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_981_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_982_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_982_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_982_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_982_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_983_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_983_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_983_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_983_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_984_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_984_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_984_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_984_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_985_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_985_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_985_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_985_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_986_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_986_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_986_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_986_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_987_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_987_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_987_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_987_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_988_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_988_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_988_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_988_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_989_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_989_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_989_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_989_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_990_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_990_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_990_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_990_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_991_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_991_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_991_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_991_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_992_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_992_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_992_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_992_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_993_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_993_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_993_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_993_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_994_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_994_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_994_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_994_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_995_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_995_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_995_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_995_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_996_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_996_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_996_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_996_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_997_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_997_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_997_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_997_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_998_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_998_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_998_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_998_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_999_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_999_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_999_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_999_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1000_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1000_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1000_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1000_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1001_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1001_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1001_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1001_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1002_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1002_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1002_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1002_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1003_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1003_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1003_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1003_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1004_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1004_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1004_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1004_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1005_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1005_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1005_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1005_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1006_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1006_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1006_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1006_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1007_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1007_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1007_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1007_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1008_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1008_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1008_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1008_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1009_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1009_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1009_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1009_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1010_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1010_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1010_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1010_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1011_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1011_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1011_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1011_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1012_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1012_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1012_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1012_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1013_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1013_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1013_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1013_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1014_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1014_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1014_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1014_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1015_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1015_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1015_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1015_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1016_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1016_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1016_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1016_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1017_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1017_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1017_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1017_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1018_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1018_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1018_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1018_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1019_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1019_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1019_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1019_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1020_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1020_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1020_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1020_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1021_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1021_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1021_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1021_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1022_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1022_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1022_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1022_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1023_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1023_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1023_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1023_en; // @[DM.scala 12:29]
  wire [31:0] RAM_MPORT_1024_data; // @[DM.scala 12:29]
  wire [9:0] RAM_MPORT_1024_addr; // @[DM.scala 12:29]
  wire  RAM_MPORT_1024_mask; // @[DM.scala 12:29]
  wire  RAM_MPORT_1024_en; // @[DM.scala 12:29]
  assign RAM_io_RD_MPORT_en = 1'h1;
  assign RAM_io_RD_MPORT_addr = io_Addr[11:2];
  assign RAM_io_RD_MPORT_data = RAM[RAM_io_RD_MPORT_addr]; // @[DM.scala 12:29]
  assign RAM_MPORT_data = 32'h0;
  assign RAM_MPORT_addr = 10'h0;
  assign RAM_MPORT_mask = 1'h1;
  assign RAM_MPORT_en = reset;
  assign RAM_MPORT_1_data = 32'h0;
  assign RAM_MPORT_1_addr = 10'h1;
  assign RAM_MPORT_1_mask = 1'h1;
  assign RAM_MPORT_1_en = reset;
  assign RAM_MPORT_2_data = 32'h0;
  assign RAM_MPORT_2_addr = 10'h2;
  assign RAM_MPORT_2_mask = 1'h1;
  assign RAM_MPORT_2_en = reset;
  assign RAM_MPORT_3_data = 32'h0;
  assign RAM_MPORT_3_addr = 10'h3;
  assign RAM_MPORT_3_mask = 1'h1;
  assign RAM_MPORT_3_en = reset;
  assign RAM_MPORT_4_data = 32'h0;
  assign RAM_MPORT_4_addr = 10'h4;
  assign RAM_MPORT_4_mask = 1'h1;
  assign RAM_MPORT_4_en = reset;
  assign RAM_MPORT_5_data = 32'h0;
  assign RAM_MPORT_5_addr = 10'h5;
  assign RAM_MPORT_5_mask = 1'h1;
  assign RAM_MPORT_5_en = reset;
  assign RAM_MPORT_6_data = 32'h0;
  assign RAM_MPORT_6_addr = 10'h6;
  assign RAM_MPORT_6_mask = 1'h1;
  assign RAM_MPORT_6_en = reset;
  assign RAM_MPORT_7_data = 32'h0;
  assign RAM_MPORT_7_addr = 10'h7;
  assign RAM_MPORT_7_mask = 1'h1;
  assign RAM_MPORT_7_en = reset;
  assign RAM_MPORT_8_data = 32'h0;
  assign RAM_MPORT_8_addr = 10'h8;
  assign RAM_MPORT_8_mask = 1'h1;
  assign RAM_MPORT_8_en = reset;
  assign RAM_MPORT_9_data = 32'h0;
  assign RAM_MPORT_9_addr = 10'h9;
  assign RAM_MPORT_9_mask = 1'h1;
  assign RAM_MPORT_9_en = reset;
  assign RAM_MPORT_10_data = 32'h0;
  assign RAM_MPORT_10_addr = 10'ha;
  assign RAM_MPORT_10_mask = 1'h1;
  assign RAM_MPORT_10_en = reset;
  assign RAM_MPORT_11_data = 32'h0;
  assign RAM_MPORT_11_addr = 10'hb;
  assign RAM_MPORT_11_mask = 1'h1;
  assign RAM_MPORT_11_en = reset;
  assign RAM_MPORT_12_data = 32'h0;
  assign RAM_MPORT_12_addr = 10'hc;
  assign RAM_MPORT_12_mask = 1'h1;
  assign RAM_MPORT_12_en = reset;
  assign RAM_MPORT_13_data = 32'h0;
  assign RAM_MPORT_13_addr = 10'hd;
  assign RAM_MPORT_13_mask = 1'h1;
  assign RAM_MPORT_13_en = reset;
  assign RAM_MPORT_14_data = 32'h0;
  assign RAM_MPORT_14_addr = 10'he;
  assign RAM_MPORT_14_mask = 1'h1;
  assign RAM_MPORT_14_en = reset;
  assign RAM_MPORT_15_data = 32'h0;
  assign RAM_MPORT_15_addr = 10'hf;
  assign RAM_MPORT_15_mask = 1'h1;
  assign RAM_MPORT_15_en = reset;
  assign RAM_MPORT_16_data = 32'h0;
  assign RAM_MPORT_16_addr = 10'h10;
  assign RAM_MPORT_16_mask = 1'h1;
  assign RAM_MPORT_16_en = reset;
  assign RAM_MPORT_17_data = 32'h0;
  assign RAM_MPORT_17_addr = 10'h11;
  assign RAM_MPORT_17_mask = 1'h1;
  assign RAM_MPORT_17_en = reset;
  assign RAM_MPORT_18_data = 32'h0;
  assign RAM_MPORT_18_addr = 10'h12;
  assign RAM_MPORT_18_mask = 1'h1;
  assign RAM_MPORT_18_en = reset;
  assign RAM_MPORT_19_data = 32'h0;
  assign RAM_MPORT_19_addr = 10'h13;
  assign RAM_MPORT_19_mask = 1'h1;
  assign RAM_MPORT_19_en = reset;
  assign RAM_MPORT_20_data = 32'h0;
  assign RAM_MPORT_20_addr = 10'h14;
  assign RAM_MPORT_20_mask = 1'h1;
  assign RAM_MPORT_20_en = reset;
  assign RAM_MPORT_21_data = 32'h0;
  assign RAM_MPORT_21_addr = 10'h15;
  assign RAM_MPORT_21_mask = 1'h1;
  assign RAM_MPORT_21_en = reset;
  assign RAM_MPORT_22_data = 32'h0;
  assign RAM_MPORT_22_addr = 10'h16;
  assign RAM_MPORT_22_mask = 1'h1;
  assign RAM_MPORT_22_en = reset;
  assign RAM_MPORT_23_data = 32'h0;
  assign RAM_MPORT_23_addr = 10'h17;
  assign RAM_MPORT_23_mask = 1'h1;
  assign RAM_MPORT_23_en = reset;
  assign RAM_MPORT_24_data = 32'h0;
  assign RAM_MPORT_24_addr = 10'h18;
  assign RAM_MPORT_24_mask = 1'h1;
  assign RAM_MPORT_24_en = reset;
  assign RAM_MPORT_25_data = 32'h0;
  assign RAM_MPORT_25_addr = 10'h19;
  assign RAM_MPORT_25_mask = 1'h1;
  assign RAM_MPORT_25_en = reset;
  assign RAM_MPORT_26_data = 32'h0;
  assign RAM_MPORT_26_addr = 10'h1a;
  assign RAM_MPORT_26_mask = 1'h1;
  assign RAM_MPORT_26_en = reset;
  assign RAM_MPORT_27_data = 32'h0;
  assign RAM_MPORT_27_addr = 10'h1b;
  assign RAM_MPORT_27_mask = 1'h1;
  assign RAM_MPORT_27_en = reset;
  assign RAM_MPORT_28_data = 32'h0;
  assign RAM_MPORT_28_addr = 10'h1c;
  assign RAM_MPORT_28_mask = 1'h1;
  assign RAM_MPORT_28_en = reset;
  assign RAM_MPORT_29_data = 32'h0;
  assign RAM_MPORT_29_addr = 10'h1d;
  assign RAM_MPORT_29_mask = 1'h1;
  assign RAM_MPORT_29_en = reset;
  assign RAM_MPORT_30_data = 32'h0;
  assign RAM_MPORT_30_addr = 10'h1e;
  assign RAM_MPORT_30_mask = 1'h1;
  assign RAM_MPORT_30_en = reset;
  assign RAM_MPORT_31_data = 32'h0;
  assign RAM_MPORT_31_addr = 10'h1f;
  assign RAM_MPORT_31_mask = 1'h1;
  assign RAM_MPORT_31_en = reset;
  assign RAM_MPORT_32_data = 32'h0;
  assign RAM_MPORT_32_addr = 10'h20;
  assign RAM_MPORT_32_mask = 1'h1;
  assign RAM_MPORT_32_en = reset;
  assign RAM_MPORT_33_data = 32'h0;
  assign RAM_MPORT_33_addr = 10'h21;
  assign RAM_MPORT_33_mask = 1'h1;
  assign RAM_MPORT_33_en = reset;
  assign RAM_MPORT_34_data = 32'h0;
  assign RAM_MPORT_34_addr = 10'h22;
  assign RAM_MPORT_34_mask = 1'h1;
  assign RAM_MPORT_34_en = reset;
  assign RAM_MPORT_35_data = 32'h0;
  assign RAM_MPORT_35_addr = 10'h23;
  assign RAM_MPORT_35_mask = 1'h1;
  assign RAM_MPORT_35_en = reset;
  assign RAM_MPORT_36_data = 32'h0;
  assign RAM_MPORT_36_addr = 10'h24;
  assign RAM_MPORT_36_mask = 1'h1;
  assign RAM_MPORT_36_en = reset;
  assign RAM_MPORT_37_data = 32'h0;
  assign RAM_MPORT_37_addr = 10'h25;
  assign RAM_MPORT_37_mask = 1'h1;
  assign RAM_MPORT_37_en = reset;
  assign RAM_MPORT_38_data = 32'h0;
  assign RAM_MPORT_38_addr = 10'h26;
  assign RAM_MPORT_38_mask = 1'h1;
  assign RAM_MPORT_38_en = reset;
  assign RAM_MPORT_39_data = 32'h0;
  assign RAM_MPORT_39_addr = 10'h27;
  assign RAM_MPORT_39_mask = 1'h1;
  assign RAM_MPORT_39_en = reset;
  assign RAM_MPORT_40_data = 32'h0;
  assign RAM_MPORT_40_addr = 10'h28;
  assign RAM_MPORT_40_mask = 1'h1;
  assign RAM_MPORT_40_en = reset;
  assign RAM_MPORT_41_data = 32'h0;
  assign RAM_MPORT_41_addr = 10'h29;
  assign RAM_MPORT_41_mask = 1'h1;
  assign RAM_MPORT_41_en = reset;
  assign RAM_MPORT_42_data = 32'h0;
  assign RAM_MPORT_42_addr = 10'h2a;
  assign RAM_MPORT_42_mask = 1'h1;
  assign RAM_MPORT_42_en = reset;
  assign RAM_MPORT_43_data = 32'h0;
  assign RAM_MPORT_43_addr = 10'h2b;
  assign RAM_MPORT_43_mask = 1'h1;
  assign RAM_MPORT_43_en = reset;
  assign RAM_MPORT_44_data = 32'h0;
  assign RAM_MPORT_44_addr = 10'h2c;
  assign RAM_MPORT_44_mask = 1'h1;
  assign RAM_MPORT_44_en = reset;
  assign RAM_MPORT_45_data = 32'h0;
  assign RAM_MPORT_45_addr = 10'h2d;
  assign RAM_MPORT_45_mask = 1'h1;
  assign RAM_MPORT_45_en = reset;
  assign RAM_MPORT_46_data = 32'h0;
  assign RAM_MPORT_46_addr = 10'h2e;
  assign RAM_MPORT_46_mask = 1'h1;
  assign RAM_MPORT_46_en = reset;
  assign RAM_MPORT_47_data = 32'h0;
  assign RAM_MPORT_47_addr = 10'h2f;
  assign RAM_MPORT_47_mask = 1'h1;
  assign RAM_MPORT_47_en = reset;
  assign RAM_MPORT_48_data = 32'h0;
  assign RAM_MPORT_48_addr = 10'h30;
  assign RAM_MPORT_48_mask = 1'h1;
  assign RAM_MPORT_48_en = reset;
  assign RAM_MPORT_49_data = 32'h0;
  assign RAM_MPORT_49_addr = 10'h31;
  assign RAM_MPORT_49_mask = 1'h1;
  assign RAM_MPORT_49_en = reset;
  assign RAM_MPORT_50_data = 32'h0;
  assign RAM_MPORT_50_addr = 10'h32;
  assign RAM_MPORT_50_mask = 1'h1;
  assign RAM_MPORT_50_en = reset;
  assign RAM_MPORT_51_data = 32'h0;
  assign RAM_MPORT_51_addr = 10'h33;
  assign RAM_MPORT_51_mask = 1'h1;
  assign RAM_MPORT_51_en = reset;
  assign RAM_MPORT_52_data = 32'h0;
  assign RAM_MPORT_52_addr = 10'h34;
  assign RAM_MPORT_52_mask = 1'h1;
  assign RAM_MPORT_52_en = reset;
  assign RAM_MPORT_53_data = 32'h0;
  assign RAM_MPORT_53_addr = 10'h35;
  assign RAM_MPORT_53_mask = 1'h1;
  assign RAM_MPORT_53_en = reset;
  assign RAM_MPORT_54_data = 32'h0;
  assign RAM_MPORT_54_addr = 10'h36;
  assign RAM_MPORT_54_mask = 1'h1;
  assign RAM_MPORT_54_en = reset;
  assign RAM_MPORT_55_data = 32'h0;
  assign RAM_MPORT_55_addr = 10'h37;
  assign RAM_MPORT_55_mask = 1'h1;
  assign RAM_MPORT_55_en = reset;
  assign RAM_MPORT_56_data = 32'h0;
  assign RAM_MPORT_56_addr = 10'h38;
  assign RAM_MPORT_56_mask = 1'h1;
  assign RAM_MPORT_56_en = reset;
  assign RAM_MPORT_57_data = 32'h0;
  assign RAM_MPORT_57_addr = 10'h39;
  assign RAM_MPORT_57_mask = 1'h1;
  assign RAM_MPORT_57_en = reset;
  assign RAM_MPORT_58_data = 32'h0;
  assign RAM_MPORT_58_addr = 10'h3a;
  assign RAM_MPORT_58_mask = 1'h1;
  assign RAM_MPORT_58_en = reset;
  assign RAM_MPORT_59_data = 32'h0;
  assign RAM_MPORT_59_addr = 10'h3b;
  assign RAM_MPORT_59_mask = 1'h1;
  assign RAM_MPORT_59_en = reset;
  assign RAM_MPORT_60_data = 32'h0;
  assign RAM_MPORT_60_addr = 10'h3c;
  assign RAM_MPORT_60_mask = 1'h1;
  assign RAM_MPORT_60_en = reset;
  assign RAM_MPORT_61_data = 32'h0;
  assign RAM_MPORT_61_addr = 10'h3d;
  assign RAM_MPORT_61_mask = 1'h1;
  assign RAM_MPORT_61_en = reset;
  assign RAM_MPORT_62_data = 32'h0;
  assign RAM_MPORT_62_addr = 10'h3e;
  assign RAM_MPORT_62_mask = 1'h1;
  assign RAM_MPORT_62_en = reset;
  assign RAM_MPORT_63_data = 32'h0;
  assign RAM_MPORT_63_addr = 10'h3f;
  assign RAM_MPORT_63_mask = 1'h1;
  assign RAM_MPORT_63_en = reset;
  assign RAM_MPORT_64_data = 32'h0;
  assign RAM_MPORT_64_addr = 10'h40;
  assign RAM_MPORT_64_mask = 1'h1;
  assign RAM_MPORT_64_en = reset;
  assign RAM_MPORT_65_data = 32'h0;
  assign RAM_MPORT_65_addr = 10'h41;
  assign RAM_MPORT_65_mask = 1'h1;
  assign RAM_MPORT_65_en = reset;
  assign RAM_MPORT_66_data = 32'h0;
  assign RAM_MPORT_66_addr = 10'h42;
  assign RAM_MPORT_66_mask = 1'h1;
  assign RAM_MPORT_66_en = reset;
  assign RAM_MPORT_67_data = 32'h0;
  assign RAM_MPORT_67_addr = 10'h43;
  assign RAM_MPORT_67_mask = 1'h1;
  assign RAM_MPORT_67_en = reset;
  assign RAM_MPORT_68_data = 32'h0;
  assign RAM_MPORT_68_addr = 10'h44;
  assign RAM_MPORT_68_mask = 1'h1;
  assign RAM_MPORT_68_en = reset;
  assign RAM_MPORT_69_data = 32'h0;
  assign RAM_MPORT_69_addr = 10'h45;
  assign RAM_MPORT_69_mask = 1'h1;
  assign RAM_MPORT_69_en = reset;
  assign RAM_MPORT_70_data = 32'h0;
  assign RAM_MPORT_70_addr = 10'h46;
  assign RAM_MPORT_70_mask = 1'h1;
  assign RAM_MPORT_70_en = reset;
  assign RAM_MPORT_71_data = 32'h0;
  assign RAM_MPORT_71_addr = 10'h47;
  assign RAM_MPORT_71_mask = 1'h1;
  assign RAM_MPORT_71_en = reset;
  assign RAM_MPORT_72_data = 32'h0;
  assign RAM_MPORT_72_addr = 10'h48;
  assign RAM_MPORT_72_mask = 1'h1;
  assign RAM_MPORT_72_en = reset;
  assign RAM_MPORT_73_data = 32'h0;
  assign RAM_MPORT_73_addr = 10'h49;
  assign RAM_MPORT_73_mask = 1'h1;
  assign RAM_MPORT_73_en = reset;
  assign RAM_MPORT_74_data = 32'h0;
  assign RAM_MPORT_74_addr = 10'h4a;
  assign RAM_MPORT_74_mask = 1'h1;
  assign RAM_MPORT_74_en = reset;
  assign RAM_MPORT_75_data = 32'h0;
  assign RAM_MPORT_75_addr = 10'h4b;
  assign RAM_MPORT_75_mask = 1'h1;
  assign RAM_MPORT_75_en = reset;
  assign RAM_MPORT_76_data = 32'h0;
  assign RAM_MPORT_76_addr = 10'h4c;
  assign RAM_MPORT_76_mask = 1'h1;
  assign RAM_MPORT_76_en = reset;
  assign RAM_MPORT_77_data = 32'h0;
  assign RAM_MPORT_77_addr = 10'h4d;
  assign RAM_MPORT_77_mask = 1'h1;
  assign RAM_MPORT_77_en = reset;
  assign RAM_MPORT_78_data = 32'h0;
  assign RAM_MPORT_78_addr = 10'h4e;
  assign RAM_MPORT_78_mask = 1'h1;
  assign RAM_MPORT_78_en = reset;
  assign RAM_MPORT_79_data = 32'h0;
  assign RAM_MPORT_79_addr = 10'h4f;
  assign RAM_MPORT_79_mask = 1'h1;
  assign RAM_MPORT_79_en = reset;
  assign RAM_MPORT_80_data = 32'h0;
  assign RAM_MPORT_80_addr = 10'h50;
  assign RAM_MPORT_80_mask = 1'h1;
  assign RAM_MPORT_80_en = reset;
  assign RAM_MPORT_81_data = 32'h0;
  assign RAM_MPORT_81_addr = 10'h51;
  assign RAM_MPORT_81_mask = 1'h1;
  assign RAM_MPORT_81_en = reset;
  assign RAM_MPORT_82_data = 32'h0;
  assign RAM_MPORT_82_addr = 10'h52;
  assign RAM_MPORT_82_mask = 1'h1;
  assign RAM_MPORT_82_en = reset;
  assign RAM_MPORT_83_data = 32'h0;
  assign RAM_MPORT_83_addr = 10'h53;
  assign RAM_MPORT_83_mask = 1'h1;
  assign RAM_MPORT_83_en = reset;
  assign RAM_MPORT_84_data = 32'h0;
  assign RAM_MPORT_84_addr = 10'h54;
  assign RAM_MPORT_84_mask = 1'h1;
  assign RAM_MPORT_84_en = reset;
  assign RAM_MPORT_85_data = 32'h0;
  assign RAM_MPORT_85_addr = 10'h55;
  assign RAM_MPORT_85_mask = 1'h1;
  assign RAM_MPORT_85_en = reset;
  assign RAM_MPORT_86_data = 32'h0;
  assign RAM_MPORT_86_addr = 10'h56;
  assign RAM_MPORT_86_mask = 1'h1;
  assign RAM_MPORT_86_en = reset;
  assign RAM_MPORT_87_data = 32'h0;
  assign RAM_MPORT_87_addr = 10'h57;
  assign RAM_MPORT_87_mask = 1'h1;
  assign RAM_MPORT_87_en = reset;
  assign RAM_MPORT_88_data = 32'h0;
  assign RAM_MPORT_88_addr = 10'h58;
  assign RAM_MPORT_88_mask = 1'h1;
  assign RAM_MPORT_88_en = reset;
  assign RAM_MPORT_89_data = 32'h0;
  assign RAM_MPORT_89_addr = 10'h59;
  assign RAM_MPORT_89_mask = 1'h1;
  assign RAM_MPORT_89_en = reset;
  assign RAM_MPORT_90_data = 32'h0;
  assign RAM_MPORT_90_addr = 10'h5a;
  assign RAM_MPORT_90_mask = 1'h1;
  assign RAM_MPORT_90_en = reset;
  assign RAM_MPORT_91_data = 32'h0;
  assign RAM_MPORT_91_addr = 10'h5b;
  assign RAM_MPORT_91_mask = 1'h1;
  assign RAM_MPORT_91_en = reset;
  assign RAM_MPORT_92_data = 32'h0;
  assign RAM_MPORT_92_addr = 10'h5c;
  assign RAM_MPORT_92_mask = 1'h1;
  assign RAM_MPORT_92_en = reset;
  assign RAM_MPORT_93_data = 32'h0;
  assign RAM_MPORT_93_addr = 10'h5d;
  assign RAM_MPORT_93_mask = 1'h1;
  assign RAM_MPORT_93_en = reset;
  assign RAM_MPORT_94_data = 32'h0;
  assign RAM_MPORT_94_addr = 10'h5e;
  assign RAM_MPORT_94_mask = 1'h1;
  assign RAM_MPORT_94_en = reset;
  assign RAM_MPORT_95_data = 32'h0;
  assign RAM_MPORT_95_addr = 10'h5f;
  assign RAM_MPORT_95_mask = 1'h1;
  assign RAM_MPORT_95_en = reset;
  assign RAM_MPORT_96_data = 32'h0;
  assign RAM_MPORT_96_addr = 10'h60;
  assign RAM_MPORT_96_mask = 1'h1;
  assign RAM_MPORT_96_en = reset;
  assign RAM_MPORT_97_data = 32'h0;
  assign RAM_MPORT_97_addr = 10'h61;
  assign RAM_MPORT_97_mask = 1'h1;
  assign RAM_MPORT_97_en = reset;
  assign RAM_MPORT_98_data = 32'h0;
  assign RAM_MPORT_98_addr = 10'h62;
  assign RAM_MPORT_98_mask = 1'h1;
  assign RAM_MPORT_98_en = reset;
  assign RAM_MPORT_99_data = 32'h0;
  assign RAM_MPORT_99_addr = 10'h63;
  assign RAM_MPORT_99_mask = 1'h1;
  assign RAM_MPORT_99_en = reset;
  assign RAM_MPORT_100_data = 32'h0;
  assign RAM_MPORT_100_addr = 10'h64;
  assign RAM_MPORT_100_mask = 1'h1;
  assign RAM_MPORT_100_en = reset;
  assign RAM_MPORT_101_data = 32'h0;
  assign RAM_MPORT_101_addr = 10'h65;
  assign RAM_MPORT_101_mask = 1'h1;
  assign RAM_MPORT_101_en = reset;
  assign RAM_MPORT_102_data = 32'h0;
  assign RAM_MPORT_102_addr = 10'h66;
  assign RAM_MPORT_102_mask = 1'h1;
  assign RAM_MPORT_102_en = reset;
  assign RAM_MPORT_103_data = 32'h0;
  assign RAM_MPORT_103_addr = 10'h67;
  assign RAM_MPORT_103_mask = 1'h1;
  assign RAM_MPORT_103_en = reset;
  assign RAM_MPORT_104_data = 32'h0;
  assign RAM_MPORT_104_addr = 10'h68;
  assign RAM_MPORT_104_mask = 1'h1;
  assign RAM_MPORT_104_en = reset;
  assign RAM_MPORT_105_data = 32'h0;
  assign RAM_MPORT_105_addr = 10'h69;
  assign RAM_MPORT_105_mask = 1'h1;
  assign RAM_MPORT_105_en = reset;
  assign RAM_MPORT_106_data = 32'h0;
  assign RAM_MPORT_106_addr = 10'h6a;
  assign RAM_MPORT_106_mask = 1'h1;
  assign RAM_MPORT_106_en = reset;
  assign RAM_MPORT_107_data = 32'h0;
  assign RAM_MPORT_107_addr = 10'h6b;
  assign RAM_MPORT_107_mask = 1'h1;
  assign RAM_MPORT_107_en = reset;
  assign RAM_MPORT_108_data = 32'h0;
  assign RAM_MPORT_108_addr = 10'h6c;
  assign RAM_MPORT_108_mask = 1'h1;
  assign RAM_MPORT_108_en = reset;
  assign RAM_MPORT_109_data = 32'h0;
  assign RAM_MPORT_109_addr = 10'h6d;
  assign RAM_MPORT_109_mask = 1'h1;
  assign RAM_MPORT_109_en = reset;
  assign RAM_MPORT_110_data = 32'h0;
  assign RAM_MPORT_110_addr = 10'h6e;
  assign RAM_MPORT_110_mask = 1'h1;
  assign RAM_MPORT_110_en = reset;
  assign RAM_MPORT_111_data = 32'h0;
  assign RAM_MPORT_111_addr = 10'h6f;
  assign RAM_MPORT_111_mask = 1'h1;
  assign RAM_MPORT_111_en = reset;
  assign RAM_MPORT_112_data = 32'h0;
  assign RAM_MPORT_112_addr = 10'h70;
  assign RAM_MPORT_112_mask = 1'h1;
  assign RAM_MPORT_112_en = reset;
  assign RAM_MPORT_113_data = 32'h0;
  assign RAM_MPORT_113_addr = 10'h71;
  assign RAM_MPORT_113_mask = 1'h1;
  assign RAM_MPORT_113_en = reset;
  assign RAM_MPORT_114_data = 32'h0;
  assign RAM_MPORT_114_addr = 10'h72;
  assign RAM_MPORT_114_mask = 1'h1;
  assign RAM_MPORT_114_en = reset;
  assign RAM_MPORT_115_data = 32'h0;
  assign RAM_MPORT_115_addr = 10'h73;
  assign RAM_MPORT_115_mask = 1'h1;
  assign RAM_MPORT_115_en = reset;
  assign RAM_MPORT_116_data = 32'h0;
  assign RAM_MPORT_116_addr = 10'h74;
  assign RAM_MPORT_116_mask = 1'h1;
  assign RAM_MPORT_116_en = reset;
  assign RAM_MPORT_117_data = 32'h0;
  assign RAM_MPORT_117_addr = 10'h75;
  assign RAM_MPORT_117_mask = 1'h1;
  assign RAM_MPORT_117_en = reset;
  assign RAM_MPORT_118_data = 32'h0;
  assign RAM_MPORT_118_addr = 10'h76;
  assign RAM_MPORT_118_mask = 1'h1;
  assign RAM_MPORT_118_en = reset;
  assign RAM_MPORT_119_data = 32'h0;
  assign RAM_MPORT_119_addr = 10'h77;
  assign RAM_MPORT_119_mask = 1'h1;
  assign RAM_MPORT_119_en = reset;
  assign RAM_MPORT_120_data = 32'h0;
  assign RAM_MPORT_120_addr = 10'h78;
  assign RAM_MPORT_120_mask = 1'h1;
  assign RAM_MPORT_120_en = reset;
  assign RAM_MPORT_121_data = 32'h0;
  assign RAM_MPORT_121_addr = 10'h79;
  assign RAM_MPORT_121_mask = 1'h1;
  assign RAM_MPORT_121_en = reset;
  assign RAM_MPORT_122_data = 32'h0;
  assign RAM_MPORT_122_addr = 10'h7a;
  assign RAM_MPORT_122_mask = 1'h1;
  assign RAM_MPORT_122_en = reset;
  assign RAM_MPORT_123_data = 32'h0;
  assign RAM_MPORT_123_addr = 10'h7b;
  assign RAM_MPORT_123_mask = 1'h1;
  assign RAM_MPORT_123_en = reset;
  assign RAM_MPORT_124_data = 32'h0;
  assign RAM_MPORT_124_addr = 10'h7c;
  assign RAM_MPORT_124_mask = 1'h1;
  assign RAM_MPORT_124_en = reset;
  assign RAM_MPORT_125_data = 32'h0;
  assign RAM_MPORT_125_addr = 10'h7d;
  assign RAM_MPORT_125_mask = 1'h1;
  assign RAM_MPORT_125_en = reset;
  assign RAM_MPORT_126_data = 32'h0;
  assign RAM_MPORT_126_addr = 10'h7e;
  assign RAM_MPORT_126_mask = 1'h1;
  assign RAM_MPORT_126_en = reset;
  assign RAM_MPORT_127_data = 32'h0;
  assign RAM_MPORT_127_addr = 10'h7f;
  assign RAM_MPORT_127_mask = 1'h1;
  assign RAM_MPORT_127_en = reset;
  assign RAM_MPORT_128_data = 32'h0;
  assign RAM_MPORT_128_addr = 10'h80;
  assign RAM_MPORT_128_mask = 1'h1;
  assign RAM_MPORT_128_en = reset;
  assign RAM_MPORT_129_data = 32'h0;
  assign RAM_MPORT_129_addr = 10'h81;
  assign RAM_MPORT_129_mask = 1'h1;
  assign RAM_MPORT_129_en = reset;
  assign RAM_MPORT_130_data = 32'h0;
  assign RAM_MPORT_130_addr = 10'h82;
  assign RAM_MPORT_130_mask = 1'h1;
  assign RAM_MPORT_130_en = reset;
  assign RAM_MPORT_131_data = 32'h0;
  assign RAM_MPORT_131_addr = 10'h83;
  assign RAM_MPORT_131_mask = 1'h1;
  assign RAM_MPORT_131_en = reset;
  assign RAM_MPORT_132_data = 32'h0;
  assign RAM_MPORT_132_addr = 10'h84;
  assign RAM_MPORT_132_mask = 1'h1;
  assign RAM_MPORT_132_en = reset;
  assign RAM_MPORT_133_data = 32'h0;
  assign RAM_MPORT_133_addr = 10'h85;
  assign RAM_MPORT_133_mask = 1'h1;
  assign RAM_MPORT_133_en = reset;
  assign RAM_MPORT_134_data = 32'h0;
  assign RAM_MPORT_134_addr = 10'h86;
  assign RAM_MPORT_134_mask = 1'h1;
  assign RAM_MPORT_134_en = reset;
  assign RAM_MPORT_135_data = 32'h0;
  assign RAM_MPORT_135_addr = 10'h87;
  assign RAM_MPORT_135_mask = 1'h1;
  assign RAM_MPORT_135_en = reset;
  assign RAM_MPORT_136_data = 32'h0;
  assign RAM_MPORT_136_addr = 10'h88;
  assign RAM_MPORT_136_mask = 1'h1;
  assign RAM_MPORT_136_en = reset;
  assign RAM_MPORT_137_data = 32'h0;
  assign RAM_MPORT_137_addr = 10'h89;
  assign RAM_MPORT_137_mask = 1'h1;
  assign RAM_MPORT_137_en = reset;
  assign RAM_MPORT_138_data = 32'h0;
  assign RAM_MPORT_138_addr = 10'h8a;
  assign RAM_MPORT_138_mask = 1'h1;
  assign RAM_MPORT_138_en = reset;
  assign RAM_MPORT_139_data = 32'h0;
  assign RAM_MPORT_139_addr = 10'h8b;
  assign RAM_MPORT_139_mask = 1'h1;
  assign RAM_MPORT_139_en = reset;
  assign RAM_MPORT_140_data = 32'h0;
  assign RAM_MPORT_140_addr = 10'h8c;
  assign RAM_MPORT_140_mask = 1'h1;
  assign RAM_MPORT_140_en = reset;
  assign RAM_MPORT_141_data = 32'h0;
  assign RAM_MPORT_141_addr = 10'h8d;
  assign RAM_MPORT_141_mask = 1'h1;
  assign RAM_MPORT_141_en = reset;
  assign RAM_MPORT_142_data = 32'h0;
  assign RAM_MPORT_142_addr = 10'h8e;
  assign RAM_MPORT_142_mask = 1'h1;
  assign RAM_MPORT_142_en = reset;
  assign RAM_MPORT_143_data = 32'h0;
  assign RAM_MPORT_143_addr = 10'h8f;
  assign RAM_MPORT_143_mask = 1'h1;
  assign RAM_MPORT_143_en = reset;
  assign RAM_MPORT_144_data = 32'h0;
  assign RAM_MPORT_144_addr = 10'h90;
  assign RAM_MPORT_144_mask = 1'h1;
  assign RAM_MPORT_144_en = reset;
  assign RAM_MPORT_145_data = 32'h0;
  assign RAM_MPORT_145_addr = 10'h91;
  assign RAM_MPORT_145_mask = 1'h1;
  assign RAM_MPORT_145_en = reset;
  assign RAM_MPORT_146_data = 32'h0;
  assign RAM_MPORT_146_addr = 10'h92;
  assign RAM_MPORT_146_mask = 1'h1;
  assign RAM_MPORT_146_en = reset;
  assign RAM_MPORT_147_data = 32'h0;
  assign RAM_MPORT_147_addr = 10'h93;
  assign RAM_MPORT_147_mask = 1'h1;
  assign RAM_MPORT_147_en = reset;
  assign RAM_MPORT_148_data = 32'h0;
  assign RAM_MPORT_148_addr = 10'h94;
  assign RAM_MPORT_148_mask = 1'h1;
  assign RAM_MPORT_148_en = reset;
  assign RAM_MPORT_149_data = 32'h0;
  assign RAM_MPORT_149_addr = 10'h95;
  assign RAM_MPORT_149_mask = 1'h1;
  assign RAM_MPORT_149_en = reset;
  assign RAM_MPORT_150_data = 32'h0;
  assign RAM_MPORT_150_addr = 10'h96;
  assign RAM_MPORT_150_mask = 1'h1;
  assign RAM_MPORT_150_en = reset;
  assign RAM_MPORT_151_data = 32'h0;
  assign RAM_MPORT_151_addr = 10'h97;
  assign RAM_MPORT_151_mask = 1'h1;
  assign RAM_MPORT_151_en = reset;
  assign RAM_MPORT_152_data = 32'h0;
  assign RAM_MPORT_152_addr = 10'h98;
  assign RAM_MPORT_152_mask = 1'h1;
  assign RAM_MPORT_152_en = reset;
  assign RAM_MPORT_153_data = 32'h0;
  assign RAM_MPORT_153_addr = 10'h99;
  assign RAM_MPORT_153_mask = 1'h1;
  assign RAM_MPORT_153_en = reset;
  assign RAM_MPORT_154_data = 32'h0;
  assign RAM_MPORT_154_addr = 10'h9a;
  assign RAM_MPORT_154_mask = 1'h1;
  assign RAM_MPORT_154_en = reset;
  assign RAM_MPORT_155_data = 32'h0;
  assign RAM_MPORT_155_addr = 10'h9b;
  assign RAM_MPORT_155_mask = 1'h1;
  assign RAM_MPORT_155_en = reset;
  assign RAM_MPORT_156_data = 32'h0;
  assign RAM_MPORT_156_addr = 10'h9c;
  assign RAM_MPORT_156_mask = 1'h1;
  assign RAM_MPORT_156_en = reset;
  assign RAM_MPORT_157_data = 32'h0;
  assign RAM_MPORT_157_addr = 10'h9d;
  assign RAM_MPORT_157_mask = 1'h1;
  assign RAM_MPORT_157_en = reset;
  assign RAM_MPORT_158_data = 32'h0;
  assign RAM_MPORT_158_addr = 10'h9e;
  assign RAM_MPORT_158_mask = 1'h1;
  assign RAM_MPORT_158_en = reset;
  assign RAM_MPORT_159_data = 32'h0;
  assign RAM_MPORT_159_addr = 10'h9f;
  assign RAM_MPORT_159_mask = 1'h1;
  assign RAM_MPORT_159_en = reset;
  assign RAM_MPORT_160_data = 32'h0;
  assign RAM_MPORT_160_addr = 10'ha0;
  assign RAM_MPORT_160_mask = 1'h1;
  assign RAM_MPORT_160_en = reset;
  assign RAM_MPORT_161_data = 32'h0;
  assign RAM_MPORT_161_addr = 10'ha1;
  assign RAM_MPORT_161_mask = 1'h1;
  assign RAM_MPORT_161_en = reset;
  assign RAM_MPORT_162_data = 32'h0;
  assign RAM_MPORT_162_addr = 10'ha2;
  assign RAM_MPORT_162_mask = 1'h1;
  assign RAM_MPORT_162_en = reset;
  assign RAM_MPORT_163_data = 32'h0;
  assign RAM_MPORT_163_addr = 10'ha3;
  assign RAM_MPORT_163_mask = 1'h1;
  assign RAM_MPORT_163_en = reset;
  assign RAM_MPORT_164_data = 32'h0;
  assign RAM_MPORT_164_addr = 10'ha4;
  assign RAM_MPORT_164_mask = 1'h1;
  assign RAM_MPORT_164_en = reset;
  assign RAM_MPORT_165_data = 32'h0;
  assign RAM_MPORT_165_addr = 10'ha5;
  assign RAM_MPORT_165_mask = 1'h1;
  assign RAM_MPORT_165_en = reset;
  assign RAM_MPORT_166_data = 32'h0;
  assign RAM_MPORT_166_addr = 10'ha6;
  assign RAM_MPORT_166_mask = 1'h1;
  assign RAM_MPORT_166_en = reset;
  assign RAM_MPORT_167_data = 32'h0;
  assign RAM_MPORT_167_addr = 10'ha7;
  assign RAM_MPORT_167_mask = 1'h1;
  assign RAM_MPORT_167_en = reset;
  assign RAM_MPORT_168_data = 32'h0;
  assign RAM_MPORT_168_addr = 10'ha8;
  assign RAM_MPORT_168_mask = 1'h1;
  assign RAM_MPORT_168_en = reset;
  assign RAM_MPORT_169_data = 32'h0;
  assign RAM_MPORT_169_addr = 10'ha9;
  assign RAM_MPORT_169_mask = 1'h1;
  assign RAM_MPORT_169_en = reset;
  assign RAM_MPORT_170_data = 32'h0;
  assign RAM_MPORT_170_addr = 10'haa;
  assign RAM_MPORT_170_mask = 1'h1;
  assign RAM_MPORT_170_en = reset;
  assign RAM_MPORT_171_data = 32'h0;
  assign RAM_MPORT_171_addr = 10'hab;
  assign RAM_MPORT_171_mask = 1'h1;
  assign RAM_MPORT_171_en = reset;
  assign RAM_MPORT_172_data = 32'h0;
  assign RAM_MPORT_172_addr = 10'hac;
  assign RAM_MPORT_172_mask = 1'h1;
  assign RAM_MPORT_172_en = reset;
  assign RAM_MPORT_173_data = 32'h0;
  assign RAM_MPORT_173_addr = 10'had;
  assign RAM_MPORT_173_mask = 1'h1;
  assign RAM_MPORT_173_en = reset;
  assign RAM_MPORT_174_data = 32'h0;
  assign RAM_MPORT_174_addr = 10'hae;
  assign RAM_MPORT_174_mask = 1'h1;
  assign RAM_MPORT_174_en = reset;
  assign RAM_MPORT_175_data = 32'h0;
  assign RAM_MPORT_175_addr = 10'haf;
  assign RAM_MPORT_175_mask = 1'h1;
  assign RAM_MPORT_175_en = reset;
  assign RAM_MPORT_176_data = 32'h0;
  assign RAM_MPORT_176_addr = 10'hb0;
  assign RAM_MPORT_176_mask = 1'h1;
  assign RAM_MPORT_176_en = reset;
  assign RAM_MPORT_177_data = 32'h0;
  assign RAM_MPORT_177_addr = 10'hb1;
  assign RAM_MPORT_177_mask = 1'h1;
  assign RAM_MPORT_177_en = reset;
  assign RAM_MPORT_178_data = 32'h0;
  assign RAM_MPORT_178_addr = 10'hb2;
  assign RAM_MPORT_178_mask = 1'h1;
  assign RAM_MPORT_178_en = reset;
  assign RAM_MPORT_179_data = 32'h0;
  assign RAM_MPORT_179_addr = 10'hb3;
  assign RAM_MPORT_179_mask = 1'h1;
  assign RAM_MPORT_179_en = reset;
  assign RAM_MPORT_180_data = 32'h0;
  assign RAM_MPORT_180_addr = 10'hb4;
  assign RAM_MPORT_180_mask = 1'h1;
  assign RAM_MPORT_180_en = reset;
  assign RAM_MPORT_181_data = 32'h0;
  assign RAM_MPORT_181_addr = 10'hb5;
  assign RAM_MPORT_181_mask = 1'h1;
  assign RAM_MPORT_181_en = reset;
  assign RAM_MPORT_182_data = 32'h0;
  assign RAM_MPORT_182_addr = 10'hb6;
  assign RAM_MPORT_182_mask = 1'h1;
  assign RAM_MPORT_182_en = reset;
  assign RAM_MPORT_183_data = 32'h0;
  assign RAM_MPORT_183_addr = 10'hb7;
  assign RAM_MPORT_183_mask = 1'h1;
  assign RAM_MPORT_183_en = reset;
  assign RAM_MPORT_184_data = 32'h0;
  assign RAM_MPORT_184_addr = 10'hb8;
  assign RAM_MPORT_184_mask = 1'h1;
  assign RAM_MPORT_184_en = reset;
  assign RAM_MPORT_185_data = 32'h0;
  assign RAM_MPORT_185_addr = 10'hb9;
  assign RAM_MPORT_185_mask = 1'h1;
  assign RAM_MPORT_185_en = reset;
  assign RAM_MPORT_186_data = 32'h0;
  assign RAM_MPORT_186_addr = 10'hba;
  assign RAM_MPORT_186_mask = 1'h1;
  assign RAM_MPORT_186_en = reset;
  assign RAM_MPORT_187_data = 32'h0;
  assign RAM_MPORT_187_addr = 10'hbb;
  assign RAM_MPORT_187_mask = 1'h1;
  assign RAM_MPORT_187_en = reset;
  assign RAM_MPORT_188_data = 32'h0;
  assign RAM_MPORT_188_addr = 10'hbc;
  assign RAM_MPORT_188_mask = 1'h1;
  assign RAM_MPORT_188_en = reset;
  assign RAM_MPORT_189_data = 32'h0;
  assign RAM_MPORT_189_addr = 10'hbd;
  assign RAM_MPORT_189_mask = 1'h1;
  assign RAM_MPORT_189_en = reset;
  assign RAM_MPORT_190_data = 32'h0;
  assign RAM_MPORT_190_addr = 10'hbe;
  assign RAM_MPORT_190_mask = 1'h1;
  assign RAM_MPORT_190_en = reset;
  assign RAM_MPORT_191_data = 32'h0;
  assign RAM_MPORT_191_addr = 10'hbf;
  assign RAM_MPORT_191_mask = 1'h1;
  assign RAM_MPORT_191_en = reset;
  assign RAM_MPORT_192_data = 32'h0;
  assign RAM_MPORT_192_addr = 10'hc0;
  assign RAM_MPORT_192_mask = 1'h1;
  assign RAM_MPORT_192_en = reset;
  assign RAM_MPORT_193_data = 32'h0;
  assign RAM_MPORT_193_addr = 10'hc1;
  assign RAM_MPORT_193_mask = 1'h1;
  assign RAM_MPORT_193_en = reset;
  assign RAM_MPORT_194_data = 32'h0;
  assign RAM_MPORT_194_addr = 10'hc2;
  assign RAM_MPORT_194_mask = 1'h1;
  assign RAM_MPORT_194_en = reset;
  assign RAM_MPORT_195_data = 32'h0;
  assign RAM_MPORT_195_addr = 10'hc3;
  assign RAM_MPORT_195_mask = 1'h1;
  assign RAM_MPORT_195_en = reset;
  assign RAM_MPORT_196_data = 32'h0;
  assign RAM_MPORT_196_addr = 10'hc4;
  assign RAM_MPORT_196_mask = 1'h1;
  assign RAM_MPORT_196_en = reset;
  assign RAM_MPORT_197_data = 32'h0;
  assign RAM_MPORT_197_addr = 10'hc5;
  assign RAM_MPORT_197_mask = 1'h1;
  assign RAM_MPORT_197_en = reset;
  assign RAM_MPORT_198_data = 32'h0;
  assign RAM_MPORT_198_addr = 10'hc6;
  assign RAM_MPORT_198_mask = 1'h1;
  assign RAM_MPORT_198_en = reset;
  assign RAM_MPORT_199_data = 32'h0;
  assign RAM_MPORT_199_addr = 10'hc7;
  assign RAM_MPORT_199_mask = 1'h1;
  assign RAM_MPORT_199_en = reset;
  assign RAM_MPORT_200_data = 32'h0;
  assign RAM_MPORT_200_addr = 10'hc8;
  assign RAM_MPORT_200_mask = 1'h1;
  assign RAM_MPORT_200_en = reset;
  assign RAM_MPORT_201_data = 32'h0;
  assign RAM_MPORT_201_addr = 10'hc9;
  assign RAM_MPORT_201_mask = 1'h1;
  assign RAM_MPORT_201_en = reset;
  assign RAM_MPORT_202_data = 32'h0;
  assign RAM_MPORT_202_addr = 10'hca;
  assign RAM_MPORT_202_mask = 1'h1;
  assign RAM_MPORT_202_en = reset;
  assign RAM_MPORT_203_data = 32'h0;
  assign RAM_MPORT_203_addr = 10'hcb;
  assign RAM_MPORT_203_mask = 1'h1;
  assign RAM_MPORT_203_en = reset;
  assign RAM_MPORT_204_data = 32'h0;
  assign RAM_MPORT_204_addr = 10'hcc;
  assign RAM_MPORT_204_mask = 1'h1;
  assign RAM_MPORT_204_en = reset;
  assign RAM_MPORT_205_data = 32'h0;
  assign RAM_MPORT_205_addr = 10'hcd;
  assign RAM_MPORT_205_mask = 1'h1;
  assign RAM_MPORT_205_en = reset;
  assign RAM_MPORT_206_data = 32'h0;
  assign RAM_MPORT_206_addr = 10'hce;
  assign RAM_MPORT_206_mask = 1'h1;
  assign RAM_MPORT_206_en = reset;
  assign RAM_MPORT_207_data = 32'h0;
  assign RAM_MPORT_207_addr = 10'hcf;
  assign RAM_MPORT_207_mask = 1'h1;
  assign RAM_MPORT_207_en = reset;
  assign RAM_MPORT_208_data = 32'h0;
  assign RAM_MPORT_208_addr = 10'hd0;
  assign RAM_MPORT_208_mask = 1'h1;
  assign RAM_MPORT_208_en = reset;
  assign RAM_MPORT_209_data = 32'h0;
  assign RAM_MPORT_209_addr = 10'hd1;
  assign RAM_MPORT_209_mask = 1'h1;
  assign RAM_MPORT_209_en = reset;
  assign RAM_MPORT_210_data = 32'h0;
  assign RAM_MPORT_210_addr = 10'hd2;
  assign RAM_MPORT_210_mask = 1'h1;
  assign RAM_MPORT_210_en = reset;
  assign RAM_MPORT_211_data = 32'h0;
  assign RAM_MPORT_211_addr = 10'hd3;
  assign RAM_MPORT_211_mask = 1'h1;
  assign RAM_MPORT_211_en = reset;
  assign RAM_MPORT_212_data = 32'h0;
  assign RAM_MPORT_212_addr = 10'hd4;
  assign RAM_MPORT_212_mask = 1'h1;
  assign RAM_MPORT_212_en = reset;
  assign RAM_MPORT_213_data = 32'h0;
  assign RAM_MPORT_213_addr = 10'hd5;
  assign RAM_MPORT_213_mask = 1'h1;
  assign RAM_MPORT_213_en = reset;
  assign RAM_MPORT_214_data = 32'h0;
  assign RAM_MPORT_214_addr = 10'hd6;
  assign RAM_MPORT_214_mask = 1'h1;
  assign RAM_MPORT_214_en = reset;
  assign RAM_MPORT_215_data = 32'h0;
  assign RAM_MPORT_215_addr = 10'hd7;
  assign RAM_MPORT_215_mask = 1'h1;
  assign RAM_MPORT_215_en = reset;
  assign RAM_MPORT_216_data = 32'h0;
  assign RAM_MPORT_216_addr = 10'hd8;
  assign RAM_MPORT_216_mask = 1'h1;
  assign RAM_MPORT_216_en = reset;
  assign RAM_MPORT_217_data = 32'h0;
  assign RAM_MPORT_217_addr = 10'hd9;
  assign RAM_MPORT_217_mask = 1'h1;
  assign RAM_MPORT_217_en = reset;
  assign RAM_MPORT_218_data = 32'h0;
  assign RAM_MPORT_218_addr = 10'hda;
  assign RAM_MPORT_218_mask = 1'h1;
  assign RAM_MPORT_218_en = reset;
  assign RAM_MPORT_219_data = 32'h0;
  assign RAM_MPORT_219_addr = 10'hdb;
  assign RAM_MPORT_219_mask = 1'h1;
  assign RAM_MPORT_219_en = reset;
  assign RAM_MPORT_220_data = 32'h0;
  assign RAM_MPORT_220_addr = 10'hdc;
  assign RAM_MPORT_220_mask = 1'h1;
  assign RAM_MPORT_220_en = reset;
  assign RAM_MPORT_221_data = 32'h0;
  assign RAM_MPORT_221_addr = 10'hdd;
  assign RAM_MPORT_221_mask = 1'h1;
  assign RAM_MPORT_221_en = reset;
  assign RAM_MPORT_222_data = 32'h0;
  assign RAM_MPORT_222_addr = 10'hde;
  assign RAM_MPORT_222_mask = 1'h1;
  assign RAM_MPORT_222_en = reset;
  assign RAM_MPORT_223_data = 32'h0;
  assign RAM_MPORT_223_addr = 10'hdf;
  assign RAM_MPORT_223_mask = 1'h1;
  assign RAM_MPORT_223_en = reset;
  assign RAM_MPORT_224_data = 32'h0;
  assign RAM_MPORT_224_addr = 10'he0;
  assign RAM_MPORT_224_mask = 1'h1;
  assign RAM_MPORT_224_en = reset;
  assign RAM_MPORT_225_data = 32'h0;
  assign RAM_MPORT_225_addr = 10'he1;
  assign RAM_MPORT_225_mask = 1'h1;
  assign RAM_MPORT_225_en = reset;
  assign RAM_MPORT_226_data = 32'h0;
  assign RAM_MPORT_226_addr = 10'he2;
  assign RAM_MPORT_226_mask = 1'h1;
  assign RAM_MPORT_226_en = reset;
  assign RAM_MPORT_227_data = 32'h0;
  assign RAM_MPORT_227_addr = 10'he3;
  assign RAM_MPORT_227_mask = 1'h1;
  assign RAM_MPORT_227_en = reset;
  assign RAM_MPORT_228_data = 32'h0;
  assign RAM_MPORT_228_addr = 10'he4;
  assign RAM_MPORT_228_mask = 1'h1;
  assign RAM_MPORT_228_en = reset;
  assign RAM_MPORT_229_data = 32'h0;
  assign RAM_MPORT_229_addr = 10'he5;
  assign RAM_MPORT_229_mask = 1'h1;
  assign RAM_MPORT_229_en = reset;
  assign RAM_MPORT_230_data = 32'h0;
  assign RAM_MPORT_230_addr = 10'he6;
  assign RAM_MPORT_230_mask = 1'h1;
  assign RAM_MPORT_230_en = reset;
  assign RAM_MPORT_231_data = 32'h0;
  assign RAM_MPORT_231_addr = 10'he7;
  assign RAM_MPORT_231_mask = 1'h1;
  assign RAM_MPORT_231_en = reset;
  assign RAM_MPORT_232_data = 32'h0;
  assign RAM_MPORT_232_addr = 10'he8;
  assign RAM_MPORT_232_mask = 1'h1;
  assign RAM_MPORT_232_en = reset;
  assign RAM_MPORT_233_data = 32'h0;
  assign RAM_MPORT_233_addr = 10'he9;
  assign RAM_MPORT_233_mask = 1'h1;
  assign RAM_MPORT_233_en = reset;
  assign RAM_MPORT_234_data = 32'h0;
  assign RAM_MPORT_234_addr = 10'hea;
  assign RAM_MPORT_234_mask = 1'h1;
  assign RAM_MPORT_234_en = reset;
  assign RAM_MPORT_235_data = 32'h0;
  assign RAM_MPORT_235_addr = 10'heb;
  assign RAM_MPORT_235_mask = 1'h1;
  assign RAM_MPORT_235_en = reset;
  assign RAM_MPORT_236_data = 32'h0;
  assign RAM_MPORT_236_addr = 10'hec;
  assign RAM_MPORT_236_mask = 1'h1;
  assign RAM_MPORT_236_en = reset;
  assign RAM_MPORT_237_data = 32'h0;
  assign RAM_MPORT_237_addr = 10'hed;
  assign RAM_MPORT_237_mask = 1'h1;
  assign RAM_MPORT_237_en = reset;
  assign RAM_MPORT_238_data = 32'h0;
  assign RAM_MPORT_238_addr = 10'hee;
  assign RAM_MPORT_238_mask = 1'h1;
  assign RAM_MPORT_238_en = reset;
  assign RAM_MPORT_239_data = 32'h0;
  assign RAM_MPORT_239_addr = 10'hef;
  assign RAM_MPORT_239_mask = 1'h1;
  assign RAM_MPORT_239_en = reset;
  assign RAM_MPORT_240_data = 32'h0;
  assign RAM_MPORT_240_addr = 10'hf0;
  assign RAM_MPORT_240_mask = 1'h1;
  assign RAM_MPORT_240_en = reset;
  assign RAM_MPORT_241_data = 32'h0;
  assign RAM_MPORT_241_addr = 10'hf1;
  assign RAM_MPORT_241_mask = 1'h1;
  assign RAM_MPORT_241_en = reset;
  assign RAM_MPORT_242_data = 32'h0;
  assign RAM_MPORT_242_addr = 10'hf2;
  assign RAM_MPORT_242_mask = 1'h1;
  assign RAM_MPORT_242_en = reset;
  assign RAM_MPORT_243_data = 32'h0;
  assign RAM_MPORT_243_addr = 10'hf3;
  assign RAM_MPORT_243_mask = 1'h1;
  assign RAM_MPORT_243_en = reset;
  assign RAM_MPORT_244_data = 32'h0;
  assign RAM_MPORT_244_addr = 10'hf4;
  assign RAM_MPORT_244_mask = 1'h1;
  assign RAM_MPORT_244_en = reset;
  assign RAM_MPORT_245_data = 32'h0;
  assign RAM_MPORT_245_addr = 10'hf5;
  assign RAM_MPORT_245_mask = 1'h1;
  assign RAM_MPORT_245_en = reset;
  assign RAM_MPORT_246_data = 32'h0;
  assign RAM_MPORT_246_addr = 10'hf6;
  assign RAM_MPORT_246_mask = 1'h1;
  assign RAM_MPORT_246_en = reset;
  assign RAM_MPORT_247_data = 32'h0;
  assign RAM_MPORT_247_addr = 10'hf7;
  assign RAM_MPORT_247_mask = 1'h1;
  assign RAM_MPORT_247_en = reset;
  assign RAM_MPORT_248_data = 32'h0;
  assign RAM_MPORT_248_addr = 10'hf8;
  assign RAM_MPORT_248_mask = 1'h1;
  assign RAM_MPORT_248_en = reset;
  assign RAM_MPORT_249_data = 32'h0;
  assign RAM_MPORT_249_addr = 10'hf9;
  assign RAM_MPORT_249_mask = 1'h1;
  assign RAM_MPORT_249_en = reset;
  assign RAM_MPORT_250_data = 32'h0;
  assign RAM_MPORT_250_addr = 10'hfa;
  assign RAM_MPORT_250_mask = 1'h1;
  assign RAM_MPORT_250_en = reset;
  assign RAM_MPORT_251_data = 32'h0;
  assign RAM_MPORT_251_addr = 10'hfb;
  assign RAM_MPORT_251_mask = 1'h1;
  assign RAM_MPORT_251_en = reset;
  assign RAM_MPORT_252_data = 32'h0;
  assign RAM_MPORT_252_addr = 10'hfc;
  assign RAM_MPORT_252_mask = 1'h1;
  assign RAM_MPORT_252_en = reset;
  assign RAM_MPORT_253_data = 32'h0;
  assign RAM_MPORT_253_addr = 10'hfd;
  assign RAM_MPORT_253_mask = 1'h1;
  assign RAM_MPORT_253_en = reset;
  assign RAM_MPORT_254_data = 32'h0;
  assign RAM_MPORT_254_addr = 10'hfe;
  assign RAM_MPORT_254_mask = 1'h1;
  assign RAM_MPORT_254_en = reset;
  assign RAM_MPORT_255_data = 32'h0;
  assign RAM_MPORT_255_addr = 10'hff;
  assign RAM_MPORT_255_mask = 1'h1;
  assign RAM_MPORT_255_en = reset;
  assign RAM_MPORT_256_data = 32'h0;
  assign RAM_MPORT_256_addr = 10'h100;
  assign RAM_MPORT_256_mask = 1'h1;
  assign RAM_MPORT_256_en = reset;
  assign RAM_MPORT_257_data = 32'h0;
  assign RAM_MPORT_257_addr = 10'h101;
  assign RAM_MPORT_257_mask = 1'h1;
  assign RAM_MPORT_257_en = reset;
  assign RAM_MPORT_258_data = 32'h0;
  assign RAM_MPORT_258_addr = 10'h102;
  assign RAM_MPORT_258_mask = 1'h1;
  assign RAM_MPORT_258_en = reset;
  assign RAM_MPORT_259_data = 32'h0;
  assign RAM_MPORT_259_addr = 10'h103;
  assign RAM_MPORT_259_mask = 1'h1;
  assign RAM_MPORT_259_en = reset;
  assign RAM_MPORT_260_data = 32'h0;
  assign RAM_MPORT_260_addr = 10'h104;
  assign RAM_MPORT_260_mask = 1'h1;
  assign RAM_MPORT_260_en = reset;
  assign RAM_MPORT_261_data = 32'h0;
  assign RAM_MPORT_261_addr = 10'h105;
  assign RAM_MPORT_261_mask = 1'h1;
  assign RAM_MPORT_261_en = reset;
  assign RAM_MPORT_262_data = 32'h0;
  assign RAM_MPORT_262_addr = 10'h106;
  assign RAM_MPORT_262_mask = 1'h1;
  assign RAM_MPORT_262_en = reset;
  assign RAM_MPORT_263_data = 32'h0;
  assign RAM_MPORT_263_addr = 10'h107;
  assign RAM_MPORT_263_mask = 1'h1;
  assign RAM_MPORT_263_en = reset;
  assign RAM_MPORT_264_data = 32'h0;
  assign RAM_MPORT_264_addr = 10'h108;
  assign RAM_MPORT_264_mask = 1'h1;
  assign RAM_MPORT_264_en = reset;
  assign RAM_MPORT_265_data = 32'h0;
  assign RAM_MPORT_265_addr = 10'h109;
  assign RAM_MPORT_265_mask = 1'h1;
  assign RAM_MPORT_265_en = reset;
  assign RAM_MPORT_266_data = 32'h0;
  assign RAM_MPORT_266_addr = 10'h10a;
  assign RAM_MPORT_266_mask = 1'h1;
  assign RAM_MPORT_266_en = reset;
  assign RAM_MPORT_267_data = 32'h0;
  assign RAM_MPORT_267_addr = 10'h10b;
  assign RAM_MPORT_267_mask = 1'h1;
  assign RAM_MPORT_267_en = reset;
  assign RAM_MPORT_268_data = 32'h0;
  assign RAM_MPORT_268_addr = 10'h10c;
  assign RAM_MPORT_268_mask = 1'h1;
  assign RAM_MPORT_268_en = reset;
  assign RAM_MPORT_269_data = 32'h0;
  assign RAM_MPORT_269_addr = 10'h10d;
  assign RAM_MPORT_269_mask = 1'h1;
  assign RAM_MPORT_269_en = reset;
  assign RAM_MPORT_270_data = 32'h0;
  assign RAM_MPORT_270_addr = 10'h10e;
  assign RAM_MPORT_270_mask = 1'h1;
  assign RAM_MPORT_270_en = reset;
  assign RAM_MPORT_271_data = 32'h0;
  assign RAM_MPORT_271_addr = 10'h10f;
  assign RAM_MPORT_271_mask = 1'h1;
  assign RAM_MPORT_271_en = reset;
  assign RAM_MPORT_272_data = 32'h0;
  assign RAM_MPORT_272_addr = 10'h110;
  assign RAM_MPORT_272_mask = 1'h1;
  assign RAM_MPORT_272_en = reset;
  assign RAM_MPORT_273_data = 32'h0;
  assign RAM_MPORT_273_addr = 10'h111;
  assign RAM_MPORT_273_mask = 1'h1;
  assign RAM_MPORT_273_en = reset;
  assign RAM_MPORT_274_data = 32'h0;
  assign RAM_MPORT_274_addr = 10'h112;
  assign RAM_MPORT_274_mask = 1'h1;
  assign RAM_MPORT_274_en = reset;
  assign RAM_MPORT_275_data = 32'h0;
  assign RAM_MPORT_275_addr = 10'h113;
  assign RAM_MPORT_275_mask = 1'h1;
  assign RAM_MPORT_275_en = reset;
  assign RAM_MPORT_276_data = 32'h0;
  assign RAM_MPORT_276_addr = 10'h114;
  assign RAM_MPORT_276_mask = 1'h1;
  assign RAM_MPORT_276_en = reset;
  assign RAM_MPORT_277_data = 32'h0;
  assign RAM_MPORT_277_addr = 10'h115;
  assign RAM_MPORT_277_mask = 1'h1;
  assign RAM_MPORT_277_en = reset;
  assign RAM_MPORT_278_data = 32'h0;
  assign RAM_MPORT_278_addr = 10'h116;
  assign RAM_MPORT_278_mask = 1'h1;
  assign RAM_MPORT_278_en = reset;
  assign RAM_MPORT_279_data = 32'h0;
  assign RAM_MPORT_279_addr = 10'h117;
  assign RAM_MPORT_279_mask = 1'h1;
  assign RAM_MPORT_279_en = reset;
  assign RAM_MPORT_280_data = 32'h0;
  assign RAM_MPORT_280_addr = 10'h118;
  assign RAM_MPORT_280_mask = 1'h1;
  assign RAM_MPORT_280_en = reset;
  assign RAM_MPORT_281_data = 32'h0;
  assign RAM_MPORT_281_addr = 10'h119;
  assign RAM_MPORT_281_mask = 1'h1;
  assign RAM_MPORT_281_en = reset;
  assign RAM_MPORT_282_data = 32'h0;
  assign RAM_MPORT_282_addr = 10'h11a;
  assign RAM_MPORT_282_mask = 1'h1;
  assign RAM_MPORT_282_en = reset;
  assign RAM_MPORT_283_data = 32'h0;
  assign RAM_MPORT_283_addr = 10'h11b;
  assign RAM_MPORT_283_mask = 1'h1;
  assign RAM_MPORT_283_en = reset;
  assign RAM_MPORT_284_data = 32'h0;
  assign RAM_MPORT_284_addr = 10'h11c;
  assign RAM_MPORT_284_mask = 1'h1;
  assign RAM_MPORT_284_en = reset;
  assign RAM_MPORT_285_data = 32'h0;
  assign RAM_MPORT_285_addr = 10'h11d;
  assign RAM_MPORT_285_mask = 1'h1;
  assign RAM_MPORT_285_en = reset;
  assign RAM_MPORT_286_data = 32'h0;
  assign RAM_MPORT_286_addr = 10'h11e;
  assign RAM_MPORT_286_mask = 1'h1;
  assign RAM_MPORT_286_en = reset;
  assign RAM_MPORT_287_data = 32'h0;
  assign RAM_MPORT_287_addr = 10'h11f;
  assign RAM_MPORT_287_mask = 1'h1;
  assign RAM_MPORT_287_en = reset;
  assign RAM_MPORT_288_data = 32'h0;
  assign RAM_MPORT_288_addr = 10'h120;
  assign RAM_MPORT_288_mask = 1'h1;
  assign RAM_MPORT_288_en = reset;
  assign RAM_MPORT_289_data = 32'h0;
  assign RAM_MPORT_289_addr = 10'h121;
  assign RAM_MPORT_289_mask = 1'h1;
  assign RAM_MPORT_289_en = reset;
  assign RAM_MPORT_290_data = 32'h0;
  assign RAM_MPORT_290_addr = 10'h122;
  assign RAM_MPORT_290_mask = 1'h1;
  assign RAM_MPORT_290_en = reset;
  assign RAM_MPORT_291_data = 32'h0;
  assign RAM_MPORT_291_addr = 10'h123;
  assign RAM_MPORT_291_mask = 1'h1;
  assign RAM_MPORT_291_en = reset;
  assign RAM_MPORT_292_data = 32'h0;
  assign RAM_MPORT_292_addr = 10'h124;
  assign RAM_MPORT_292_mask = 1'h1;
  assign RAM_MPORT_292_en = reset;
  assign RAM_MPORT_293_data = 32'h0;
  assign RAM_MPORT_293_addr = 10'h125;
  assign RAM_MPORT_293_mask = 1'h1;
  assign RAM_MPORT_293_en = reset;
  assign RAM_MPORT_294_data = 32'h0;
  assign RAM_MPORT_294_addr = 10'h126;
  assign RAM_MPORT_294_mask = 1'h1;
  assign RAM_MPORT_294_en = reset;
  assign RAM_MPORT_295_data = 32'h0;
  assign RAM_MPORT_295_addr = 10'h127;
  assign RAM_MPORT_295_mask = 1'h1;
  assign RAM_MPORT_295_en = reset;
  assign RAM_MPORT_296_data = 32'h0;
  assign RAM_MPORT_296_addr = 10'h128;
  assign RAM_MPORT_296_mask = 1'h1;
  assign RAM_MPORT_296_en = reset;
  assign RAM_MPORT_297_data = 32'h0;
  assign RAM_MPORT_297_addr = 10'h129;
  assign RAM_MPORT_297_mask = 1'h1;
  assign RAM_MPORT_297_en = reset;
  assign RAM_MPORT_298_data = 32'h0;
  assign RAM_MPORT_298_addr = 10'h12a;
  assign RAM_MPORT_298_mask = 1'h1;
  assign RAM_MPORT_298_en = reset;
  assign RAM_MPORT_299_data = 32'h0;
  assign RAM_MPORT_299_addr = 10'h12b;
  assign RAM_MPORT_299_mask = 1'h1;
  assign RAM_MPORT_299_en = reset;
  assign RAM_MPORT_300_data = 32'h0;
  assign RAM_MPORT_300_addr = 10'h12c;
  assign RAM_MPORT_300_mask = 1'h1;
  assign RAM_MPORT_300_en = reset;
  assign RAM_MPORT_301_data = 32'h0;
  assign RAM_MPORT_301_addr = 10'h12d;
  assign RAM_MPORT_301_mask = 1'h1;
  assign RAM_MPORT_301_en = reset;
  assign RAM_MPORT_302_data = 32'h0;
  assign RAM_MPORT_302_addr = 10'h12e;
  assign RAM_MPORT_302_mask = 1'h1;
  assign RAM_MPORT_302_en = reset;
  assign RAM_MPORT_303_data = 32'h0;
  assign RAM_MPORT_303_addr = 10'h12f;
  assign RAM_MPORT_303_mask = 1'h1;
  assign RAM_MPORT_303_en = reset;
  assign RAM_MPORT_304_data = 32'h0;
  assign RAM_MPORT_304_addr = 10'h130;
  assign RAM_MPORT_304_mask = 1'h1;
  assign RAM_MPORT_304_en = reset;
  assign RAM_MPORT_305_data = 32'h0;
  assign RAM_MPORT_305_addr = 10'h131;
  assign RAM_MPORT_305_mask = 1'h1;
  assign RAM_MPORT_305_en = reset;
  assign RAM_MPORT_306_data = 32'h0;
  assign RAM_MPORT_306_addr = 10'h132;
  assign RAM_MPORT_306_mask = 1'h1;
  assign RAM_MPORT_306_en = reset;
  assign RAM_MPORT_307_data = 32'h0;
  assign RAM_MPORT_307_addr = 10'h133;
  assign RAM_MPORT_307_mask = 1'h1;
  assign RAM_MPORT_307_en = reset;
  assign RAM_MPORT_308_data = 32'h0;
  assign RAM_MPORT_308_addr = 10'h134;
  assign RAM_MPORT_308_mask = 1'h1;
  assign RAM_MPORT_308_en = reset;
  assign RAM_MPORT_309_data = 32'h0;
  assign RAM_MPORT_309_addr = 10'h135;
  assign RAM_MPORT_309_mask = 1'h1;
  assign RAM_MPORT_309_en = reset;
  assign RAM_MPORT_310_data = 32'h0;
  assign RAM_MPORT_310_addr = 10'h136;
  assign RAM_MPORT_310_mask = 1'h1;
  assign RAM_MPORT_310_en = reset;
  assign RAM_MPORT_311_data = 32'h0;
  assign RAM_MPORT_311_addr = 10'h137;
  assign RAM_MPORT_311_mask = 1'h1;
  assign RAM_MPORT_311_en = reset;
  assign RAM_MPORT_312_data = 32'h0;
  assign RAM_MPORT_312_addr = 10'h138;
  assign RAM_MPORT_312_mask = 1'h1;
  assign RAM_MPORT_312_en = reset;
  assign RAM_MPORT_313_data = 32'h0;
  assign RAM_MPORT_313_addr = 10'h139;
  assign RAM_MPORT_313_mask = 1'h1;
  assign RAM_MPORT_313_en = reset;
  assign RAM_MPORT_314_data = 32'h0;
  assign RAM_MPORT_314_addr = 10'h13a;
  assign RAM_MPORT_314_mask = 1'h1;
  assign RAM_MPORT_314_en = reset;
  assign RAM_MPORT_315_data = 32'h0;
  assign RAM_MPORT_315_addr = 10'h13b;
  assign RAM_MPORT_315_mask = 1'h1;
  assign RAM_MPORT_315_en = reset;
  assign RAM_MPORT_316_data = 32'h0;
  assign RAM_MPORT_316_addr = 10'h13c;
  assign RAM_MPORT_316_mask = 1'h1;
  assign RAM_MPORT_316_en = reset;
  assign RAM_MPORT_317_data = 32'h0;
  assign RAM_MPORT_317_addr = 10'h13d;
  assign RAM_MPORT_317_mask = 1'h1;
  assign RAM_MPORT_317_en = reset;
  assign RAM_MPORT_318_data = 32'h0;
  assign RAM_MPORT_318_addr = 10'h13e;
  assign RAM_MPORT_318_mask = 1'h1;
  assign RAM_MPORT_318_en = reset;
  assign RAM_MPORT_319_data = 32'h0;
  assign RAM_MPORT_319_addr = 10'h13f;
  assign RAM_MPORT_319_mask = 1'h1;
  assign RAM_MPORT_319_en = reset;
  assign RAM_MPORT_320_data = 32'h0;
  assign RAM_MPORT_320_addr = 10'h140;
  assign RAM_MPORT_320_mask = 1'h1;
  assign RAM_MPORT_320_en = reset;
  assign RAM_MPORT_321_data = 32'h0;
  assign RAM_MPORT_321_addr = 10'h141;
  assign RAM_MPORT_321_mask = 1'h1;
  assign RAM_MPORT_321_en = reset;
  assign RAM_MPORT_322_data = 32'h0;
  assign RAM_MPORT_322_addr = 10'h142;
  assign RAM_MPORT_322_mask = 1'h1;
  assign RAM_MPORT_322_en = reset;
  assign RAM_MPORT_323_data = 32'h0;
  assign RAM_MPORT_323_addr = 10'h143;
  assign RAM_MPORT_323_mask = 1'h1;
  assign RAM_MPORT_323_en = reset;
  assign RAM_MPORT_324_data = 32'h0;
  assign RAM_MPORT_324_addr = 10'h144;
  assign RAM_MPORT_324_mask = 1'h1;
  assign RAM_MPORT_324_en = reset;
  assign RAM_MPORT_325_data = 32'h0;
  assign RAM_MPORT_325_addr = 10'h145;
  assign RAM_MPORT_325_mask = 1'h1;
  assign RAM_MPORT_325_en = reset;
  assign RAM_MPORT_326_data = 32'h0;
  assign RAM_MPORT_326_addr = 10'h146;
  assign RAM_MPORT_326_mask = 1'h1;
  assign RAM_MPORT_326_en = reset;
  assign RAM_MPORT_327_data = 32'h0;
  assign RAM_MPORT_327_addr = 10'h147;
  assign RAM_MPORT_327_mask = 1'h1;
  assign RAM_MPORT_327_en = reset;
  assign RAM_MPORT_328_data = 32'h0;
  assign RAM_MPORT_328_addr = 10'h148;
  assign RAM_MPORT_328_mask = 1'h1;
  assign RAM_MPORT_328_en = reset;
  assign RAM_MPORT_329_data = 32'h0;
  assign RAM_MPORT_329_addr = 10'h149;
  assign RAM_MPORT_329_mask = 1'h1;
  assign RAM_MPORT_329_en = reset;
  assign RAM_MPORT_330_data = 32'h0;
  assign RAM_MPORT_330_addr = 10'h14a;
  assign RAM_MPORT_330_mask = 1'h1;
  assign RAM_MPORT_330_en = reset;
  assign RAM_MPORT_331_data = 32'h0;
  assign RAM_MPORT_331_addr = 10'h14b;
  assign RAM_MPORT_331_mask = 1'h1;
  assign RAM_MPORT_331_en = reset;
  assign RAM_MPORT_332_data = 32'h0;
  assign RAM_MPORT_332_addr = 10'h14c;
  assign RAM_MPORT_332_mask = 1'h1;
  assign RAM_MPORT_332_en = reset;
  assign RAM_MPORT_333_data = 32'h0;
  assign RAM_MPORT_333_addr = 10'h14d;
  assign RAM_MPORT_333_mask = 1'h1;
  assign RAM_MPORT_333_en = reset;
  assign RAM_MPORT_334_data = 32'h0;
  assign RAM_MPORT_334_addr = 10'h14e;
  assign RAM_MPORT_334_mask = 1'h1;
  assign RAM_MPORT_334_en = reset;
  assign RAM_MPORT_335_data = 32'h0;
  assign RAM_MPORT_335_addr = 10'h14f;
  assign RAM_MPORT_335_mask = 1'h1;
  assign RAM_MPORT_335_en = reset;
  assign RAM_MPORT_336_data = 32'h0;
  assign RAM_MPORT_336_addr = 10'h150;
  assign RAM_MPORT_336_mask = 1'h1;
  assign RAM_MPORT_336_en = reset;
  assign RAM_MPORT_337_data = 32'h0;
  assign RAM_MPORT_337_addr = 10'h151;
  assign RAM_MPORT_337_mask = 1'h1;
  assign RAM_MPORT_337_en = reset;
  assign RAM_MPORT_338_data = 32'h0;
  assign RAM_MPORT_338_addr = 10'h152;
  assign RAM_MPORT_338_mask = 1'h1;
  assign RAM_MPORT_338_en = reset;
  assign RAM_MPORT_339_data = 32'h0;
  assign RAM_MPORT_339_addr = 10'h153;
  assign RAM_MPORT_339_mask = 1'h1;
  assign RAM_MPORT_339_en = reset;
  assign RAM_MPORT_340_data = 32'h0;
  assign RAM_MPORT_340_addr = 10'h154;
  assign RAM_MPORT_340_mask = 1'h1;
  assign RAM_MPORT_340_en = reset;
  assign RAM_MPORT_341_data = 32'h0;
  assign RAM_MPORT_341_addr = 10'h155;
  assign RAM_MPORT_341_mask = 1'h1;
  assign RAM_MPORT_341_en = reset;
  assign RAM_MPORT_342_data = 32'h0;
  assign RAM_MPORT_342_addr = 10'h156;
  assign RAM_MPORT_342_mask = 1'h1;
  assign RAM_MPORT_342_en = reset;
  assign RAM_MPORT_343_data = 32'h0;
  assign RAM_MPORT_343_addr = 10'h157;
  assign RAM_MPORT_343_mask = 1'h1;
  assign RAM_MPORT_343_en = reset;
  assign RAM_MPORT_344_data = 32'h0;
  assign RAM_MPORT_344_addr = 10'h158;
  assign RAM_MPORT_344_mask = 1'h1;
  assign RAM_MPORT_344_en = reset;
  assign RAM_MPORT_345_data = 32'h0;
  assign RAM_MPORT_345_addr = 10'h159;
  assign RAM_MPORT_345_mask = 1'h1;
  assign RAM_MPORT_345_en = reset;
  assign RAM_MPORT_346_data = 32'h0;
  assign RAM_MPORT_346_addr = 10'h15a;
  assign RAM_MPORT_346_mask = 1'h1;
  assign RAM_MPORT_346_en = reset;
  assign RAM_MPORT_347_data = 32'h0;
  assign RAM_MPORT_347_addr = 10'h15b;
  assign RAM_MPORT_347_mask = 1'h1;
  assign RAM_MPORT_347_en = reset;
  assign RAM_MPORT_348_data = 32'h0;
  assign RAM_MPORT_348_addr = 10'h15c;
  assign RAM_MPORT_348_mask = 1'h1;
  assign RAM_MPORT_348_en = reset;
  assign RAM_MPORT_349_data = 32'h0;
  assign RAM_MPORT_349_addr = 10'h15d;
  assign RAM_MPORT_349_mask = 1'h1;
  assign RAM_MPORT_349_en = reset;
  assign RAM_MPORT_350_data = 32'h0;
  assign RAM_MPORT_350_addr = 10'h15e;
  assign RAM_MPORT_350_mask = 1'h1;
  assign RAM_MPORT_350_en = reset;
  assign RAM_MPORT_351_data = 32'h0;
  assign RAM_MPORT_351_addr = 10'h15f;
  assign RAM_MPORT_351_mask = 1'h1;
  assign RAM_MPORT_351_en = reset;
  assign RAM_MPORT_352_data = 32'h0;
  assign RAM_MPORT_352_addr = 10'h160;
  assign RAM_MPORT_352_mask = 1'h1;
  assign RAM_MPORT_352_en = reset;
  assign RAM_MPORT_353_data = 32'h0;
  assign RAM_MPORT_353_addr = 10'h161;
  assign RAM_MPORT_353_mask = 1'h1;
  assign RAM_MPORT_353_en = reset;
  assign RAM_MPORT_354_data = 32'h0;
  assign RAM_MPORT_354_addr = 10'h162;
  assign RAM_MPORT_354_mask = 1'h1;
  assign RAM_MPORT_354_en = reset;
  assign RAM_MPORT_355_data = 32'h0;
  assign RAM_MPORT_355_addr = 10'h163;
  assign RAM_MPORT_355_mask = 1'h1;
  assign RAM_MPORT_355_en = reset;
  assign RAM_MPORT_356_data = 32'h0;
  assign RAM_MPORT_356_addr = 10'h164;
  assign RAM_MPORT_356_mask = 1'h1;
  assign RAM_MPORT_356_en = reset;
  assign RAM_MPORT_357_data = 32'h0;
  assign RAM_MPORT_357_addr = 10'h165;
  assign RAM_MPORT_357_mask = 1'h1;
  assign RAM_MPORT_357_en = reset;
  assign RAM_MPORT_358_data = 32'h0;
  assign RAM_MPORT_358_addr = 10'h166;
  assign RAM_MPORT_358_mask = 1'h1;
  assign RAM_MPORT_358_en = reset;
  assign RAM_MPORT_359_data = 32'h0;
  assign RAM_MPORT_359_addr = 10'h167;
  assign RAM_MPORT_359_mask = 1'h1;
  assign RAM_MPORT_359_en = reset;
  assign RAM_MPORT_360_data = 32'h0;
  assign RAM_MPORT_360_addr = 10'h168;
  assign RAM_MPORT_360_mask = 1'h1;
  assign RAM_MPORT_360_en = reset;
  assign RAM_MPORT_361_data = 32'h0;
  assign RAM_MPORT_361_addr = 10'h169;
  assign RAM_MPORT_361_mask = 1'h1;
  assign RAM_MPORT_361_en = reset;
  assign RAM_MPORT_362_data = 32'h0;
  assign RAM_MPORT_362_addr = 10'h16a;
  assign RAM_MPORT_362_mask = 1'h1;
  assign RAM_MPORT_362_en = reset;
  assign RAM_MPORT_363_data = 32'h0;
  assign RAM_MPORT_363_addr = 10'h16b;
  assign RAM_MPORT_363_mask = 1'h1;
  assign RAM_MPORT_363_en = reset;
  assign RAM_MPORT_364_data = 32'h0;
  assign RAM_MPORT_364_addr = 10'h16c;
  assign RAM_MPORT_364_mask = 1'h1;
  assign RAM_MPORT_364_en = reset;
  assign RAM_MPORT_365_data = 32'h0;
  assign RAM_MPORT_365_addr = 10'h16d;
  assign RAM_MPORT_365_mask = 1'h1;
  assign RAM_MPORT_365_en = reset;
  assign RAM_MPORT_366_data = 32'h0;
  assign RAM_MPORT_366_addr = 10'h16e;
  assign RAM_MPORT_366_mask = 1'h1;
  assign RAM_MPORT_366_en = reset;
  assign RAM_MPORT_367_data = 32'h0;
  assign RAM_MPORT_367_addr = 10'h16f;
  assign RAM_MPORT_367_mask = 1'h1;
  assign RAM_MPORT_367_en = reset;
  assign RAM_MPORT_368_data = 32'h0;
  assign RAM_MPORT_368_addr = 10'h170;
  assign RAM_MPORT_368_mask = 1'h1;
  assign RAM_MPORT_368_en = reset;
  assign RAM_MPORT_369_data = 32'h0;
  assign RAM_MPORT_369_addr = 10'h171;
  assign RAM_MPORT_369_mask = 1'h1;
  assign RAM_MPORT_369_en = reset;
  assign RAM_MPORT_370_data = 32'h0;
  assign RAM_MPORT_370_addr = 10'h172;
  assign RAM_MPORT_370_mask = 1'h1;
  assign RAM_MPORT_370_en = reset;
  assign RAM_MPORT_371_data = 32'h0;
  assign RAM_MPORT_371_addr = 10'h173;
  assign RAM_MPORT_371_mask = 1'h1;
  assign RAM_MPORT_371_en = reset;
  assign RAM_MPORT_372_data = 32'h0;
  assign RAM_MPORT_372_addr = 10'h174;
  assign RAM_MPORT_372_mask = 1'h1;
  assign RAM_MPORT_372_en = reset;
  assign RAM_MPORT_373_data = 32'h0;
  assign RAM_MPORT_373_addr = 10'h175;
  assign RAM_MPORT_373_mask = 1'h1;
  assign RAM_MPORT_373_en = reset;
  assign RAM_MPORT_374_data = 32'h0;
  assign RAM_MPORT_374_addr = 10'h176;
  assign RAM_MPORT_374_mask = 1'h1;
  assign RAM_MPORT_374_en = reset;
  assign RAM_MPORT_375_data = 32'h0;
  assign RAM_MPORT_375_addr = 10'h177;
  assign RAM_MPORT_375_mask = 1'h1;
  assign RAM_MPORT_375_en = reset;
  assign RAM_MPORT_376_data = 32'h0;
  assign RAM_MPORT_376_addr = 10'h178;
  assign RAM_MPORT_376_mask = 1'h1;
  assign RAM_MPORT_376_en = reset;
  assign RAM_MPORT_377_data = 32'h0;
  assign RAM_MPORT_377_addr = 10'h179;
  assign RAM_MPORT_377_mask = 1'h1;
  assign RAM_MPORT_377_en = reset;
  assign RAM_MPORT_378_data = 32'h0;
  assign RAM_MPORT_378_addr = 10'h17a;
  assign RAM_MPORT_378_mask = 1'h1;
  assign RAM_MPORT_378_en = reset;
  assign RAM_MPORT_379_data = 32'h0;
  assign RAM_MPORT_379_addr = 10'h17b;
  assign RAM_MPORT_379_mask = 1'h1;
  assign RAM_MPORT_379_en = reset;
  assign RAM_MPORT_380_data = 32'h0;
  assign RAM_MPORT_380_addr = 10'h17c;
  assign RAM_MPORT_380_mask = 1'h1;
  assign RAM_MPORT_380_en = reset;
  assign RAM_MPORT_381_data = 32'h0;
  assign RAM_MPORT_381_addr = 10'h17d;
  assign RAM_MPORT_381_mask = 1'h1;
  assign RAM_MPORT_381_en = reset;
  assign RAM_MPORT_382_data = 32'h0;
  assign RAM_MPORT_382_addr = 10'h17e;
  assign RAM_MPORT_382_mask = 1'h1;
  assign RAM_MPORT_382_en = reset;
  assign RAM_MPORT_383_data = 32'h0;
  assign RAM_MPORT_383_addr = 10'h17f;
  assign RAM_MPORT_383_mask = 1'h1;
  assign RAM_MPORT_383_en = reset;
  assign RAM_MPORT_384_data = 32'h0;
  assign RAM_MPORT_384_addr = 10'h180;
  assign RAM_MPORT_384_mask = 1'h1;
  assign RAM_MPORT_384_en = reset;
  assign RAM_MPORT_385_data = 32'h0;
  assign RAM_MPORT_385_addr = 10'h181;
  assign RAM_MPORT_385_mask = 1'h1;
  assign RAM_MPORT_385_en = reset;
  assign RAM_MPORT_386_data = 32'h0;
  assign RAM_MPORT_386_addr = 10'h182;
  assign RAM_MPORT_386_mask = 1'h1;
  assign RAM_MPORT_386_en = reset;
  assign RAM_MPORT_387_data = 32'h0;
  assign RAM_MPORT_387_addr = 10'h183;
  assign RAM_MPORT_387_mask = 1'h1;
  assign RAM_MPORT_387_en = reset;
  assign RAM_MPORT_388_data = 32'h0;
  assign RAM_MPORT_388_addr = 10'h184;
  assign RAM_MPORT_388_mask = 1'h1;
  assign RAM_MPORT_388_en = reset;
  assign RAM_MPORT_389_data = 32'h0;
  assign RAM_MPORT_389_addr = 10'h185;
  assign RAM_MPORT_389_mask = 1'h1;
  assign RAM_MPORT_389_en = reset;
  assign RAM_MPORT_390_data = 32'h0;
  assign RAM_MPORT_390_addr = 10'h186;
  assign RAM_MPORT_390_mask = 1'h1;
  assign RAM_MPORT_390_en = reset;
  assign RAM_MPORT_391_data = 32'h0;
  assign RAM_MPORT_391_addr = 10'h187;
  assign RAM_MPORT_391_mask = 1'h1;
  assign RAM_MPORT_391_en = reset;
  assign RAM_MPORT_392_data = 32'h0;
  assign RAM_MPORT_392_addr = 10'h188;
  assign RAM_MPORT_392_mask = 1'h1;
  assign RAM_MPORT_392_en = reset;
  assign RAM_MPORT_393_data = 32'h0;
  assign RAM_MPORT_393_addr = 10'h189;
  assign RAM_MPORT_393_mask = 1'h1;
  assign RAM_MPORT_393_en = reset;
  assign RAM_MPORT_394_data = 32'h0;
  assign RAM_MPORT_394_addr = 10'h18a;
  assign RAM_MPORT_394_mask = 1'h1;
  assign RAM_MPORT_394_en = reset;
  assign RAM_MPORT_395_data = 32'h0;
  assign RAM_MPORT_395_addr = 10'h18b;
  assign RAM_MPORT_395_mask = 1'h1;
  assign RAM_MPORT_395_en = reset;
  assign RAM_MPORT_396_data = 32'h0;
  assign RAM_MPORT_396_addr = 10'h18c;
  assign RAM_MPORT_396_mask = 1'h1;
  assign RAM_MPORT_396_en = reset;
  assign RAM_MPORT_397_data = 32'h0;
  assign RAM_MPORT_397_addr = 10'h18d;
  assign RAM_MPORT_397_mask = 1'h1;
  assign RAM_MPORT_397_en = reset;
  assign RAM_MPORT_398_data = 32'h0;
  assign RAM_MPORT_398_addr = 10'h18e;
  assign RAM_MPORT_398_mask = 1'h1;
  assign RAM_MPORT_398_en = reset;
  assign RAM_MPORT_399_data = 32'h0;
  assign RAM_MPORT_399_addr = 10'h18f;
  assign RAM_MPORT_399_mask = 1'h1;
  assign RAM_MPORT_399_en = reset;
  assign RAM_MPORT_400_data = 32'h0;
  assign RAM_MPORT_400_addr = 10'h190;
  assign RAM_MPORT_400_mask = 1'h1;
  assign RAM_MPORT_400_en = reset;
  assign RAM_MPORT_401_data = 32'h0;
  assign RAM_MPORT_401_addr = 10'h191;
  assign RAM_MPORT_401_mask = 1'h1;
  assign RAM_MPORT_401_en = reset;
  assign RAM_MPORT_402_data = 32'h0;
  assign RAM_MPORT_402_addr = 10'h192;
  assign RAM_MPORT_402_mask = 1'h1;
  assign RAM_MPORT_402_en = reset;
  assign RAM_MPORT_403_data = 32'h0;
  assign RAM_MPORT_403_addr = 10'h193;
  assign RAM_MPORT_403_mask = 1'h1;
  assign RAM_MPORT_403_en = reset;
  assign RAM_MPORT_404_data = 32'h0;
  assign RAM_MPORT_404_addr = 10'h194;
  assign RAM_MPORT_404_mask = 1'h1;
  assign RAM_MPORT_404_en = reset;
  assign RAM_MPORT_405_data = 32'h0;
  assign RAM_MPORT_405_addr = 10'h195;
  assign RAM_MPORT_405_mask = 1'h1;
  assign RAM_MPORT_405_en = reset;
  assign RAM_MPORT_406_data = 32'h0;
  assign RAM_MPORT_406_addr = 10'h196;
  assign RAM_MPORT_406_mask = 1'h1;
  assign RAM_MPORT_406_en = reset;
  assign RAM_MPORT_407_data = 32'h0;
  assign RAM_MPORT_407_addr = 10'h197;
  assign RAM_MPORT_407_mask = 1'h1;
  assign RAM_MPORT_407_en = reset;
  assign RAM_MPORT_408_data = 32'h0;
  assign RAM_MPORT_408_addr = 10'h198;
  assign RAM_MPORT_408_mask = 1'h1;
  assign RAM_MPORT_408_en = reset;
  assign RAM_MPORT_409_data = 32'h0;
  assign RAM_MPORT_409_addr = 10'h199;
  assign RAM_MPORT_409_mask = 1'h1;
  assign RAM_MPORT_409_en = reset;
  assign RAM_MPORT_410_data = 32'h0;
  assign RAM_MPORT_410_addr = 10'h19a;
  assign RAM_MPORT_410_mask = 1'h1;
  assign RAM_MPORT_410_en = reset;
  assign RAM_MPORT_411_data = 32'h0;
  assign RAM_MPORT_411_addr = 10'h19b;
  assign RAM_MPORT_411_mask = 1'h1;
  assign RAM_MPORT_411_en = reset;
  assign RAM_MPORT_412_data = 32'h0;
  assign RAM_MPORT_412_addr = 10'h19c;
  assign RAM_MPORT_412_mask = 1'h1;
  assign RAM_MPORT_412_en = reset;
  assign RAM_MPORT_413_data = 32'h0;
  assign RAM_MPORT_413_addr = 10'h19d;
  assign RAM_MPORT_413_mask = 1'h1;
  assign RAM_MPORT_413_en = reset;
  assign RAM_MPORT_414_data = 32'h0;
  assign RAM_MPORT_414_addr = 10'h19e;
  assign RAM_MPORT_414_mask = 1'h1;
  assign RAM_MPORT_414_en = reset;
  assign RAM_MPORT_415_data = 32'h0;
  assign RAM_MPORT_415_addr = 10'h19f;
  assign RAM_MPORT_415_mask = 1'h1;
  assign RAM_MPORT_415_en = reset;
  assign RAM_MPORT_416_data = 32'h0;
  assign RAM_MPORT_416_addr = 10'h1a0;
  assign RAM_MPORT_416_mask = 1'h1;
  assign RAM_MPORT_416_en = reset;
  assign RAM_MPORT_417_data = 32'h0;
  assign RAM_MPORT_417_addr = 10'h1a1;
  assign RAM_MPORT_417_mask = 1'h1;
  assign RAM_MPORT_417_en = reset;
  assign RAM_MPORT_418_data = 32'h0;
  assign RAM_MPORT_418_addr = 10'h1a2;
  assign RAM_MPORT_418_mask = 1'h1;
  assign RAM_MPORT_418_en = reset;
  assign RAM_MPORT_419_data = 32'h0;
  assign RAM_MPORT_419_addr = 10'h1a3;
  assign RAM_MPORT_419_mask = 1'h1;
  assign RAM_MPORT_419_en = reset;
  assign RAM_MPORT_420_data = 32'h0;
  assign RAM_MPORT_420_addr = 10'h1a4;
  assign RAM_MPORT_420_mask = 1'h1;
  assign RAM_MPORT_420_en = reset;
  assign RAM_MPORT_421_data = 32'h0;
  assign RAM_MPORT_421_addr = 10'h1a5;
  assign RAM_MPORT_421_mask = 1'h1;
  assign RAM_MPORT_421_en = reset;
  assign RAM_MPORT_422_data = 32'h0;
  assign RAM_MPORT_422_addr = 10'h1a6;
  assign RAM_MPORT_422_mask = 1'h1;
  assign RAM_MPORT_422_en = reset;
  assign RAM_MPORT_423_data = 32'h0;
  assign RAM_MPORT_423_addr = 10'h1a7;
  assign RAM_MPORT_423_mask = 1'h1;
  assign RAM_MPORT_423_en = reset;
  assign RAM_MPORT_424_data = 32'h0;
  assign RAM_MPORT_424_addr = 10'h1a8;
  assign RAM_MPORT_424_mask = 1'h1;
  assign RAM_MPORT_424_en = reset;
  assign RAM_MPORT_425_data = 32'h0;
  assign RAM_MPORT_425_addr = 10'h1a9;
  assign RAM_MPORT_425_mask = 1'h1;
  assign RAM_MPORT_425_en = reset;
  assign RAM_MPORT_426_data = 32'h0;
  assign RAM_MPORT_426_addr = 10'h1aa;
  assign RAM_MPORT_426_mask = 1'h1;
  assign RAM_MPORT_426_en = reset;
  assign RAM_MPORT_427_data = 32'h0;
  assign RAM_MPORT_427_addr = 10'h1ab;
  assign RAM_MPORT_427_mask = 1'h1;
  assign RAM_MPORT_427_en = reset;
  assign RAM_MPORT_428_data = 32'h0;
  assign RAM_MPORT_428_addr = 10'h1ac;
  assign RAM_MPORT_428_mask = 1'h1;
  assign RAM_MPORT_428_en = reset;
  assign RAM_MPORT_429_data = 32'h0;
  assign RAM_MPORT_429_addr = 10'h1ad;
  assign RAM_MPORT_429_mask = 1'h1;
  assign RAM_MPORT_429_en = reset;
  assign RAM_MPORT_430_data = 32'h0;
  assign RAM_MPORT_430_addr = 10'h1ae;
  assign RAM_MPORT_430_mask = 1'h1;
  assign RAM_MPORT_430_en = reset;
  assign RAM_MPORT_431_data = 32'h0;
  assign RAM_MPORT_431_addr = 10'h1af;
  assign RAM_MPORT_431_mask = 1'h1;
  assign RAM_MPORT_431_en = reset;
  assign RAM_MPORT_432_data = 32'h0;
  assign RAM_MPORT_432_addr = 10'h1b0;
  assign RAM_MPORT_432_mask = 1'h1;
  assign RAM_MPORT_432_en = reset;
  assign RAM_MPORT_433_data = 32'h0;
  assign RAM_MPORT_433_addr = 10'h1b1;
  assign RAM_MPORT_433_mask = 1'h1;
  assign RAM_MPORT_433_en = reset;
  assign RAM_MPORT_434_data = 32'h0;
  assign RAM_MPORT_434_addr = 10'h1b2;
  assign RAM_MPORT_434_mask = 1'h1;
  assign RAM_MPORT_434_en = reset;
  assign RAM_MPORT_435_data = 32'h0;
  assign RAM_MPORT_435_addr = 10'h1b3;
  assign RAM_MPORT_435_mask = 1'h1;
  assign RAM_MPORT_435_en = reset;
  assign RAM_MPORT_436_data = 32'h0;
  assign RAM_MPORT_436_addr = 10'h1b4;
  assign RAM_MPORT_436_mask = 1'h1;
  assign RAM_MPORT_436_en = reset;
  assign RAM_MPORT_437_data = 32'h0;
  assign RAM_MPORT_437_addr = 10'h1b5;
  assign RAM_MPORT_437_mask = 1'h1;
  assign RAM_MPORT_437_en = reset;
  assign RAM_MPORT_438_data = 32'h0;
  assign RAM_MPORT_438_addr = 10'h1b6;
  assign RAM_MPORT_438_mask = 1'h1;
  assign RAM_MPORT_438_en = reset;
  assign RAM_MPORT_439_data = 32'h0;
  assign RAM_MPORT_439_addr = 10'h1b7;
  assign RAM_MPORT_439_mask = 1'h1;
  assign RAM_MPORT_439_en = reset;
  assign RAM_MPORT_440_data = 32'h0;
  assign RAM_MPORT_440_addr = 10'h1b8;
  assign RAM_MPORT_440_mask = 1'h1;
  assign RAM_MPORT_440_en = reset;
  assign RAM_MPORT_441_data = 32'h0;
  assign RAM_MPORT_441_addr = 10'h1b9;
  assign RAM_MPORT_441_mask = 1'h1;
  assign RAM_MPORT_441_en = reset;
  assign RAM_MPORT_442_data = 32'h0;
  assign RAM_MPORT_442_addr = 10'h1ba;
  assign RAM_MPORT_442_mask = 1'h1;
  assign RAM_MPORT_442_en = reset;
  assign RAM_MPORT_443_data = 32'h0;
  assign RAM_MPORT_443_addr = 10'h1bb;
  assign RAM_MPORT_443_mask = 1'h1;
  assign RAM_MPORT_443_en = reset;
  assign RAM_MPORT_444_data = 32'h0;
  assign RAM_MPORT_444_addr = 10'h1bc;
  assign RAM_MPORT_444_mask = 1'h1;
  assign RAM_MPORT_444_en = reset;
  assign RAM_MPORT_445_data = 32'h0;
  assign RAM_MPORT_445_addr = 10'h1bd;
  assign RAM_MPORT_445_mask = 1'h1;
  assign RAM_MPORT_445_en = reset;
  assign RAM_MPORT_446_data = 32'h0;
  assign RAM_MPORT_446_addr = 10'h1be;
  assign RAM_MPORT_446_mask = 1'h1;
  assign RAM_MPORT_446_en = reset;
  assign RAM_MPORT_447_data = 32'h0;
  assign RAM_MPORT_447_addr = 10'h1bf;
  assign RAM_MPORT_447_mask = 1'h1;
  assign RAM_MPORT_447_en = reset;
  assign RAM_MPORT_448_data = 32'h0;
  assign RAM_MPORT_448_addr = 10'h1c0;
  assign RAM_MPORT_448_mask = 1'h1;
  assign RAM_MPORT_448_en = reset;
  assign RAM_MPORT_449_data = 32'h0;
  assign RAM_MPORT_449_addr = 10'h1c1;
  assign RAM_MPORT_449_mask = 1'h1;
  assign RAM_MPORT_449_en = reset;
  assign RAM_MPORT_450_data = 32'h0;
  assign RAM_MPORT_450_addr = 10'h1c2;
  assign RAM_MPORT_450_mask = 1'h1;
  assign RAM_MPORT_450_en = reset;
  assign RAM_MPORT_451_data = 32'h0;
  assign RAM_MPORT_451_addr = 10'h1c3;
  assign RAM_MPORT_451_mask = 1'h1;
  assign RAM_MPORT_451_en = reset;
  assign RAM_MPORT_452_data = 32'h0;
  assign RAM_MPORT_452_addr = 10'h1c4;
  assign RAM_MPORT_452_mask = 1'h1;
  assign RAM_MPORT_452_en = reset;
  assign RAM_MPORT_453_data = 32'h0;
  assign RAM_MPORT_453_addr = 10'h1c5;
  assign RAM_MPORT_453_mask = 1'h1;
  assign RAM_MPORT_453_en = reset;
  assign RAM_MPORT_454_data = 32'h0;
  assign RAM_MPORT_454_addr = 10'h1c6;
  assign RAM_MPORT_454_mask = 1'h1;
  assign RAM_MPORT_454_en = reset;
  assign RAM_MPORT_455_data = 32'h0;
  assign RAM_MPORT_455_addr = 10'h1c7;
  assign RAM_MPORT_455_mask = 1'h1;
  assign RAM_MPORT_455_en = reset;
  assign RAM_MPORT_456_data = 32'h0;
  assign RAM_MPORT_456_addr = 10'h1c8;
  assign RAM_MPORT_456_mask = 1'h1;
  assign RAM_MPORT_456_en = reset;
  assign RAM_MPORT_457_data = 32'h0;
  assign RAM_MPORT_457_addr = 10'h1c9;
  assign RAM_MPORT_457_mask = 1'h1;
  assign RAM_MPORT_457_en = reset;
  assign RAM_MPORT_458_data = 32'h0;
  assign RAM_MPORT_458_addr = 10'h1ca;
  assign RAM_MPORT_458_mask = 1'h1;
  assign RAM_MPORT_458_en = reset;
  assign RAM_MPORT_459_data = 32'h0;
  assign RAM_MPORT_459_addr = 10'h1cb;
  assign RAM_MPORT_459_mask = 1'h1;
  assign RAM_MPORT_459_en = reset;
  assign RAM_MPORT_460_data = 32'h0;
  assign RAM_MPORT_460_addr = 10'h1cc;
  assign RAM_MPORT_460_mask = 1'h1;
  assign RAM_MPORT_460_en = reset;
  assign RAM_MPORT_461_data = 32'h0;
  assign RAM_MPORT_461_addr = 10'h1cd;
  assign RAM_MPORT_461_mask = 1'h1;
  assign RAM_MPORT_461_en = reset;
  assign RAM_MPORT_462_data = 32'h0;
  assign RAM_MPORT_462_addr = 10'h1ce;
  assign RAM_MPORT_462_mask = 1'h1;
  assign RAM_MPORT_462_en = reset;
  assign RAM_MPORT_463_data = 32'h0;
  assign RAM_MPORT_463_addr = 10'h1cf;
  assign RAM_MPORT_463_mask = 1'h1;
  assign RAM_MPORT_463_en = reset;
  assign RAM_MPORT_464_data = 32'h0;
  assign RAM_MPORT_464_addr = 10'h1d0;
  assign RAM_MPORT_464_mask = 1'h1;
  assign RAM_MPORT_464_en = reset;
  assign RAM_MPORT_465_data = 32'h0;
  assign RAM_MPORT_465_addr = 10'h1d1;
  assign RAM_MPORT_465_mask = 1'h1;
  assign RAM_MPORT_465_en = reset;
  assign RAM_MPORT_466_data = 32'h0;
  assign RAM_MPORT_466_addr = 10'h1d2;
  assign RAM_MPORT_466_mask = 1'h1;
  assign RAM_MPORT_466_en = reset;
  assign RAM_MPORT_467_data = 32'h0;
  assign RAM_MPORT_467_addr = 10'h1d3;
  assign RAM_MPORT_467_mask = 1'h1;
  assign RAM_MPORT_467_en = reset;
  assign RAM_MPORT_468_data = 32'h0;
  assign RAM_MPORT_468_addr = 10'h1d4;
  assign RAM_MPORT_468_mask = 1'h1;
  assign RAM_MPORT_468_en = reset;
  assign RAM_MPORT_469_data = 32'h0;
  assign RAM_MPORT_469_addr = 10'h1d5;
  assign RAM_MPORT_469_mask = 1'h1;
  assign RAM_MPORT_469_en = reset;
  assign RAM_MPORT_470_data = 32'h0;
  assign RAM_MPORT_470_addr = 10'h1d6;
  assign RAM_MPORT_470_mask = 1'h1;
  assign RAM_MPORT_470_en = reset;
  assign RAM_MPORT_471_data = 32'h0;
  assign RAM_MPORT_471_addr = 10'h1d7;
  assign RAM_MPORT_471_mask = 1'h1;
  assign RAM_MPORT_471_en = reset;
  assign RAM_MPORT_472_data = 32'h0;
  assign RAM_MPORT_472_addr = 10'h1d8;
  assign RAM_MPORT_472_mask = 1'h1;
  assign RAM_MPORT_472_en = reset;
  assign RAM_MPORT_473_data = 32'h0;
  assign RAM_MPORT_473_addr = 10'h1d9;
  assign RAM_MPORT_473_mask = 1'h1;
  assign RAM_MPORT_473_en = reset;
  assign RAM_MPORT_474_data = 32'h0;
  assign RAM_MPORT_474_addr = 10'h1da;
  assign RAM_MPORT_474_mask = 1'h1;
  assign RAM_MPORT_474_en = reset;
  assign RAM_MPORT_475_data = 32'h0;
  assign RAM_MPORT_475_addr = 10'h1db;
  assign RAM_MPORT_475_mask = 1'h1;
  assign RAM_MPORT_475_en = reset;
  assign RAM_MPORT_476_data = 32'h0;
  assign RAM_MPORT_476_addr = 10'h1dc;
  assign RAM_MPORT_476_mask = 1'h1;
  assign RAM_MPORT_476_en = reset;
  assign RAM_MPORT_477_data = 32'h0;
  assign RAM_MPORT_477_addr = 10'h1dd;
  assign RAM_MPORT_477_mask = 1'h1;
  assign RAM_MPORT_477_en = reset;
  assign RAM_MPORT_478_data = 32'h0;
  assign RAM_MPORT_478_addr = 10'h1de;
  assign RAM_MPORT_478_mask = 1'h1;
  assign RAM_MPORT_478_en = reset;
  assign RAM_MPORT_479_data = 32'h0;
  assign RAM_MPORT_479_addr = 10'h1df;
  assign RAM_MPORT_479_mask = 1'h1;
  assign RAM_MPORT_479_en = reset;
  assign RAM_MPORT_480_data = 32'h0;
  assign RAM_MPORT_480_addr = 10'h1e0;
  assign RAM_MPORT_480_mask = 1'h1;
  assign RAM_MPORT_480_en = reset;
  assign RAM_MPORT_481_data = 32'h0;
  assign RAM_MPORT_481_addr = 10'h1e1;
  assign RAM_MPORT_481_mask = 1'h1;
  assign RAM_MPORT_481_en = reset;
  assign RAM_MPORT_482_data = 32'h0;
  assign RAM_MPORT_482_addr = 10'h1e2;
  assign RAM_MPORT_482_mask = 1'h1;
  assign RAM_MPORT_482_en = reset;
  assign RAM_MPORT_483_data = 32'h0;
  assign RAM_MPORT_483_addr = 10'h1e3;
  assign RAM_MPORT_483_mask = 1'h1;
  assign RAM_MPORT_483_en = reset;
  assign RAM_MPORT_484_data = 32'h0;
  assign RAM_MPORT_484_addr = 10'h1e4;
  assign RAM_MPORT_484_mask = 1'h1;
  assign RAM_MPORT_484_en = reset;
  assign RAM_MPORT_485_data = 32'h0;
  assign RAM_MPORT_485_addr = 10'h1e5;
  assign RAM_MPORT_485_mask = 1'h1;
  assign RAM_MPORT_485_en = reset;
  assign RAM_MPORT_486_data = 32'h0;
  assign RAM_MPORT_486_addr = 10'h1e6;
  assign RAM_MPORT_486_mask = 1'h1;
  assign RAM_MPORT_486_en = reset;
  assign RAM_MPORT_487_data = 32'h0;
  assign RAM_MPORT_487_addr = 10'h1e7;
  assign RAM_MPORT_487_mask = 1'h1;
  assign RAM_MPORT_487_en = reset;
  assign RAM_MPORT_488_data = 32'h0;
  assign RAM_MPORT_488_addr = 10'h1e8;
  assign RAM_MPORT_488_mask = 1'h1;
  assign RAM_MPORT_488_en = reset;
  assign RAM_MPORT_489_data = 32'h0;
  assign RAM_MPORT_489_addr = 10'h1e9;
  assign RAM_MPORT_489_mask = 1'h1;
  assign RAM_MPORT_489_en = reset;
  assign RAM_MPORT_490_data = 32'h0;
  assign RAM_MPORT_490_addr = 10'h1ea;
  assign RAM_MPORT_490_mask = 1'h1;
  assign RAM_MPORT_490_en = reset;
  assign RAM_MPORT_491_data = 32'h0;
  assign RAM_MPORT_491_addr = 10'h1eb;
  assign RAM_MPORT_491_mask = 1'h1;
  assign RAM_MPORT_491_en = reset;
  assign RAM_MPORT_492_data = 32'h0;
  assign RAM_MPORT_492_addr = 10'h1ec;
  assign RAM_MPORT_492_mask = 1'h1;
  assign RAM_MPORT_492_en = reset;
  assign RAM_MPORT_493_data = 32'h0;
  assign RAM_MPORT_493_addr = 10'h1ed;
  assign RAM_MPORT_493_mask = 1'h1;
  assign RAM_MPORT_493_en = reset;
  assign RAM_MPORT_494_data = 32'h0;
  assign RAM_MPORT_494_addr = 10'h1ee;
  assign RAM_MPORT_494_mask = 1'h1;
  assign RAM_MPORT_494_en = reset;
  assign RAM_MPORT_495_data = 32'h0;
  assign RAM_MPORT_495_addr = 10'h1ef;
  assign RAM_MPORT_495_mask = 1'h1;
  assign RAM_MPORT_495_en = reset;
  assign RAM_MPORT_496_data = 32'h0;
  assign RAM_MPORT_496_addr = 10'h1f0;
  assign RAM_MPORT_496_mask = 1'h1;
  assign RAM_MPORT_496_en = reset;
  assign RAM_MPORT_497_data = 32'h0;
  assign RAM_MPORT_497_addr = 10'h1f1;
  assign RAM_MPORT_497_mask = 1'h1;
  assign RAM_MPORT_497_en = reset;
  assign RAM_MPORT_498_data = 32'h0;
  assign RAM_MPORT_498_addr = 10'h1f2;
  assign RAM_MPORT_498_mask = 1'h1;
  assign RAM_MPORT_498_en = reset;
  assign RAM_MPORT_499_data = 32'h0;
  assign RAM_MPORT_499_addr = 10'h1f3;
  assign RAM_MPORT_499_mask = 1'h1;
  assign RAM_MPORT_499_en = reset;
  assign RAM_MPORT_500_data = 32'h0;
  assign RAM_MPORT_500_addr = 10'h1f4;
  assign RAM_MPORT_500_mask = 1'h1;
  assign RAM_MPORT_500_en = reset;
  assign RAM_MPORT_501_data = 32'h0;
  assign RAM_MPORT_501_addr = 10'h1f5;
  assign RAM_MPORT_501_mask = 1'h1;
  assign RAM_MPORT_501_en = reset;
  assign RAM_MPORT_502_data = 32'h0;
  assign RAM_MPORT_502_addr = 10'h1f6;
  assign RAM_MPORT_502_mask = 1'h1;
  assign RAM_MPORT_502_en = reset;
  assign RAM_MPORT_503_data = 32'h0;
  assign RAM_MPORT_503_addr = 10'h1f7;
  assign RAM_MPORT_503_mask = 1'h1;
  assign RAM_MPORT_503_en = reset;
  assign RAM_MPORT_504_data = 32'h0;
  assign RAM_MPORT_504_addr = 10'h1f8;
  assign RAM_MPORT_504_mask = 1'h1;
  assign RAM_MPORT_504_en = reset;
  assign RAM_MPORT_505_data = 32'h0;
  assign RAM_MPORT_505_addr = 10'h1f9;
  assign RAM_MPORT_505_mask = 1'h1;
  assign RAM_MPORT_505_en = reset;
  assign RAM_MPORT_506_data = 32'h0;
  assign RAM_MPORT_506_addr = 10'h1fa;
  assign RAM_MPORT_506_mask = 1'h1;
  assign RAM_MPORT_506_en = reset;
  assign RAM_MPORT_507_data = 32'h0;
  assign RAM_MPORT_507_addr = 10'h1fb;
  assign RAM_MPORT_507_mask = 1'h1;
  assign RAM_MPORT_507_en = reset;
  assign RAM_MPORT_508_data = 32'h0;
  assign RAM_MPORT_508_addr = 10'h1fc;
  assign RAM_MPORT_508_mask = 1'h1;
  assign RAM_MPORT_508_en = reset;
  assign RAM_MPORT_509_data = 32'h0;
  assign RAM_MPORT_509_addr = 10'h1fd;
  assign RAM_MPORT_509_mask = 1'h1;
  assign RAM_MPORT_509_en = reset;
  assign RAM_MPORT_510_data = 32'h0;
  assign RAM_MPORT_510_addr = 10'h1fe;
  assign RAM_MPORT_510_mask = 1'h1;
  assign RAM_MPORT_510_en = reset;
  assign RAM_MPORT_511_data = 32'h0;
  assign RAM_MPORT_511_addr = 10'h1ff;
  assign RAM_MPORT_511_mask = 1'h1;
  assign RAM_MPORT_511_en = reset;
  assign RAM_MPORT_512_data = 32'h0;
  assign RAM_MPORT_512_addr = 10'h200;
  assign RAM_MPORT_512_mask = 1'h1;
  assign RAM_MPORT_512_en = reset;
  assign RAM_MPORT_513_data = 32'h0;
  assign RAM_MPORT_513_addr = 10'h201;
  assign RAM_MPORT_513_mask = 1'h1;
  assign RAM_MPORT_513_en = reset;
  assign RAM_MPORT_514_data = 32'h0;
  assign RAM_MPORT_514_addr = 10'h202;
  assign RAM_MPORT_514_mask = 1'h1;
  assign RAM_MPORT_514_en = reset;
  assign RAM_MPORT_515_data = 32'h0;
  assign RAM_MPORT_515_addr = 10'h203;
  assign RAM_MPORT_515_mask = 1'h1;
  assign RAM_MPORT_515_en = reset;
  assign RAM_MPORT_516_data = 32'h0;
  assign RAM_MPORT_516_addr = 10'h204;
  assign RAM_MPORT_516_mask = 1'h1;
  assign RAM_MPORT_516_en = reset;
  assign RAM_MPORT_517_data = 32'h0;
  assign RAM_MPORT_517_addr = 10'h205;
  assign RAM_MPORT_517_mask = 1'h1;
  assign RAM_MPORT_517_en = reset;
  assign RAM_MPORT_518_data = 32'h0;
  assign RAM_MPORT_518_addr = 10'h206;
  assign RAM_MPORT_518_mask = 1'h1;
  assign RAM_MPORT_518_en = reset;
  assign RAM_MPORT_519_data = 32'h0;
  assign RAM_MPORT_519_addr = 10'h207;
  assign RAM_MPORT_519_mask = 1'h1;
  assign RAM_MPORT_519_en = reset;
  assign RAM_MPORT_520_data = 32'h0;
  assign RAM_MPORT_520_addr = 10'h208;
  assign RAM_MPORT_520_mask = 1'h1;
  assign RAM_MPORT_520_en = reset;
  assign RAM_MPORT_521_data = 32'h0;
  assign RAM_MPORT_521_addr = 10'h209;
  assign RAM_MPORT_521_mask = 1'h1;
  assign RAM_MPORT_521_en = reset;
  assign RAM_MPORT_522_data = 32'h0;
  assign RAM_MPORT_522_addr = 10'h20a;
  assign RAM_MPORT_522_mask = 1'h1;
  assign RAM_MPORT_522_en = reset;
  assign RAM_MPORT_523_data = 32'h0;
  assign RAM_MPORT_523_addr = 10'h20b;
  assign RAM_MPORT_523_mask = 1'h1;
  assign RAM_MPORT_523_en = reset;
  assign RAM_MPORT_524_data = 32'h0;
  assign RAM_MPORT_524_addr = 10'h20c;
  assign RAM_MPORT_524_mask = 1'h1;
  assign RAM_MPORT_524_en = reset;
  assign RAM_MPORT_525_data = 32'h0;
  assign RAM_MPORT_525_addr = 10'h20d;
  assign RAM_MPORT_525_mask = 1'h1;
  assign RAM_MPORT_525_en = reset;
  assign RAM_MPORT_526_data = 32'h0;
  assign RAM_MPORT_526_addr = 10'h20e;
  assign RAM_MPORT_526_mask = 1'h1;
  assign RAM_MPORT_526_en = reset;
  assign RAM_MPORT_527_data = 32'h0;
  assign RAM_MPORT_527_addr = 10'h20f;
  assign RAM_MPORT_527_mask = 1'h1;
  assign RAM_MPORT_527_en = reset;
  assign RAM_MPORT_528_data = 32'h0;
  assign RAM_MPORT_528_addr = 10'h210;
  assign RAM_MPORT_528_mask = 1'h1;
  assign RAM_MPORT_528_en = reset;
  assign RAM_MPORT_529_data = 32'h0;
  assign RAM_MPORT_529_addr = 10'h211;
  assign RAM_MPORT_529_mask = 1'h1;
  assign RAM_MPORT_529_en = reset;
  assign RAM_MPORT_530_data = 32'h0;
  assign RAM_MPORT_530_addr = 10'h212;
  assign RAM_MPORT_530_mask = 1'h1;
  assign RAM_MPORT_530_en = reset;
  assign RAM_MPORT_531_data = 32'h0;
  assign RAM_MPORT_531_addr = 10'h213;
  assign RAM_MPORT_531_mask = 1'h1;
  assign RAM_MPORT_531_en = reset;
  assign RAM_MPORT_532_data = 32'h0;
  assign RAM_MPORT_532_addr = 10'h214;
  assign RAM_MPORT_532_mask = 1'h1;
  assign RAM_MPORT_532_en = reset;
  assign RAM_MPORT_533_data = 32'h0;
  assign RAM_MPORT_533_addr = 10'h215;
  assign RAM_MPORT_533_mask = 1'h1;
  assign RAM_MPORT_533_en = reset;
  assign RAM_MPORT_534_data = 32'h0;
  assign RAM_MPORT_534_addr = 10'h216;
  assign RAM_MPORT_534_mask = 1'h1;
  assign RAM_MPORT_534_en = reset;
  assign RAM_MPORT_535_data = 32'h0;
  assign RAM_MPORT_535_addr = 10'h217;
  assign RAM_MPORT_535_mask = 1'h1;
  assign RAM_MPORT_535_en = reset;
  assign RAM_MPORT_536_data = 32'h0;
  assign RAM_MPORT_536_addr = 10'h218;
  assign RAM_MPORT_536_mask = 1'h1;
  assign RAM_MPORT_536_en = reset;
  assign RAM_MPORT_537_data = 32'h0;
  assign RAM_MPORT_537_addr = 10'h219;
  assign RAM_MPORT_537_mask = 1'h1;
  assign RAM_MPORT_537_en = reset;
  assign RAM_MPORT_538_data = 32'h0;
  assign RAM_MPORT_538_addr = 10'h21a;
  assign RAM_MPORT_538_mask = 1'h1;
  assign RAM_MPORT_538_en = reset;
  assign RAM_MPORT_539_data = 32'h0;
  assign RAM_MPORT_539_addr = 10'h21b;
  assign RAM_MPORT_539_mask = 1'h1;
  assign RAM_MPORT_539_en = reset;
  assign RAM_MPORT_540_data = 32'h0;
  assign RAM_MPORT_540_addr = 10'h21c;
  assign RAM_MPORT_540_mask = 1'h1;
  assign RAM_MPORT_540_en = reset;
  assign RAM_MPORT_541_data = 32'h0;
  assign RAM_MPORT_541_addr = 10'h21d;
  assign RAM_MPORT_541_mask = 1'h1;
  assign RAM_MPORT_541_en = reset;
  assign RAM_MPORT_542_data = 32'h0;
  assign RAM_MPORT_542_addr = 10'h21e;
  assign RAM_MPORT_542_mask = 1'h1;
  assign RAM_MPORT_542_en = reset;
  assign RAM_MPORT_543_data = 32'h0;
  assign RAM_MPORT_543_addr = 10'h21f;
  assign RAM_MPORT_543_mask = 1'h1;
  assign RAM_MPORT_543_en = reset;
  assign RAM_MPORT_544_data = 32'h0;
  assign RAM_MPORT_544_addr = 10'h220;
  assign RAM_MPORT_544_mask = 1'h1;
  assign RAM_MPORT_544_en = reset;
  assign RAM_MPORT_545_data = 32'h0;
  assign RAM_MPORT_545_addr = 10'h221;
  assign RAM_MPORT_545_mask = 1'h1;
  assign RAM_MPORT_545_en = reset;
  assign RAM_MPORT_546_data = 32'h0;
  assign RAM_MPORT_546_addr = 10'h222;
  assign RAM_MPORT_546_mask = 1'h1;
  assign RAM_MPORT_546_en = reset;
  assign RAM_MPORT_547_data = 32'h0;
  assign RAM_MPORT_547_addr = 10'h223;
  assign RAM_MPORT_547_mask = 1'h1;
  assign RAM_MPORT_547_en = reset;
  assign RAM_MPORT_548_data = 32'h0;
  assign RAM_MPORT_548_addr = 10'h224;
  assign RAM_MPORT_548_mask = 1'h1;
  assign RAM_MPORT_548_en = reset;
  assign RAM_MPORT_549_data = 32'h0;
  assign RAM_MPORT_549_addr = 10'h225;
  assign RAM_MPORT_549_mask = 1'h1;
  assign RAM_MPORT_549_en = reset;
  assign RAM_MPORT_550_data = 32'h0;
  assign RAM_MPORT_550_addr = 10'h226;
  assign RAM_MPORT_550_mask = 1'h1;
  assign RAM_MPORT_550_en = reset;
  assign RAM_MPORT_551_data = 32'h0;
  assign RAM_MPORT_551_addr = 10'h227;
  assign RAM_MPORT_551_mask = 1'h1;
  assign RAM_MPORT_551_en = reset;
  assign RAM_MPORT_552_data = 32'h0;
  assign RAM_MPORT_552_addr = 10'h228;
  assign RAM_MPORT_552_mask = 1'h1;
  assign RAM_MPORT_552_en = reset;
  assign RAM_MPORT_553_data = 32'h0;
  assign RAM_MPORT_553_addr = 10'h229;
  assign RAM_MPORT_553_mask = 1'h1;
  assign RAM_MPORT_553_en = reset;
  assign RAM_MPORT_554_data = 32'h0;
  assign RAM_MPORT_554_addr = 10'h22a;
  assign RAM_MPORT_554_mask = 1'h1;
  assign RAM_MPORT_554_en = reset;
  assign RAM_MPORT_555_data = 32'h0;
  assign RAM_MPORT_555_addr = 10'h22b;
  assign RAM_MPORT_555_mask = 1'h1;
  assign RAM_MPORT_555_en = reset;
  assign RAM_MPORT_556_data = 32'h0;
  assign RAM_MPORT_556_addr = 10'h22c;
  assign RAM_MPORT_556_mask = 1'h1;
  assign RAM_MPORT_556_en = reset;
  assign RAM_MPORT_557_data = 32'h0;
  assign RAM_MPORT_557_addr = 10'h22d;
  assign RAM_MPORT_557_mask = 1'h1;
  assign RAM_MPORT_557_en = reset;
  assign RAM_MPORT_558_data = 32'h0;
  assign RAM_MPORT_558_addr = 10'h22e;
  assign RAM_MPORT_558_mask = 1'h1;
  assign RAM_MPORT_558_en = reset;
  assign RAM_MPORT_559_data = 32'h0;
  assign RAM_MPORT_559_addr = 10'h22f;
  assign RAM_MPORT_559_mask = 1'h1;
  assign RAM_MPORT_559_en = reset;
  assign RAM_MPORT_560_data = 32'h0;
  assign RAM_MPORT_560_addr = 10'h230;
  assign RAM_MPORT_560_mask = 1'h1;
  assign RAM_MPORT_560_en = reset;
  assign RAM_MPORT_561_data = 32'h0;
  assign RAM_MPORT_561_addr = 10'h231;
  assign RAM_MPORT_561_mask = 1'h1;
  assign RAM_MPORT_561_en = reset;
  assign RAM_MPORT_562_data = 32'h0;
  assign RAM_MPORT_562_addr = 10'h232;
  assign RAM_MPORT_562_mask = 1'h1;
  assign RAM_MPORT_562_en = reset;
  assign RAM_MPORT_563_data = 32'h0;
  assign RAM_MPORT_563_addr = 10'h233;
  assign RAM_MPORT_563_mask = 1'h1;
  assign RAM_MPORT_563_en = reset;
  assign RAM_MPORT_564_data = 32'h0;
  assign RAM_MPORT_564_addr = 10'h234;
  assign RAM_MPORT_564_mask = 1'h1;
  assign RAM_MPORT_564_en = reset;
  assign RAM_MPORT_565_data = 32'h0;
  assign RAM_MPORT_565_addr = 10'h235;
  assign RAM_MPORT_565_mask = 1'h1;
  assign RAM_MPORT_565_en = reset;
  assign RAM_MPORT_566_data = 32'h0;
  assign RAM_MPORT_566_addr = 10'h236;
  assign RAM_MPORT_566_mask = 1'h1;
  assign RAM_MPORT_566_en = reset;
  assign RAM_MPORT_567_data = 32'h0;
  assign RAM_MPORT_567_addr = 10'h237;
  assign RAM_MPORT_567_mask = 1'h1;
  assign RAM_MPORT_567_en = reset;
  assign RAM_MPORT_568_data = 32'h0;
  assign RAM_MPORT_568_addr = 10'h238;
  assign RAM_MPORT_568_mask = 1'h1;
  assign RAM_MPORT_568_en = reset;
  assign RAM_MPORT_569_data = 32'h0;
  assign RAM_MPORT_569_addr = 10'h239;
  assign RAM_MPORT_569_mask = 1'h1;
  assign RAM_MPORT_569_en = reset;
  assign RAM_MPORT_570_data = 32'h0;
  assign RAM_MPORT_570_addr = 10'h23a;
  assign RAM_MPORT_570_mask = 1'h1;
  assign RAM_MPORT_570_en = reset;
  assign RAM_MPORT_571_data = 32'h0;
  assign RAM_MPORT_571_addr = 10'h23b;
  assign RAM_MPORT_571_mask = 1'h1;
  assign RAM_MPORT_571_en = reset;
  assign RAM_MPORT_572_data = 32'h0;
  assign RAM_MPORT_572_addr = 10'h23c;
  assign RAM_MPORT_572_mask = 1'h1;
  assign RAM_MPORT_572_en = reset;
  assign RAM_MPORT_573_data = 32'h0;
  assign RAM_MPORT_573_addr = 10'h23d;
  assign RAM_MPORT_573_mask = 1'h1;
  assign RAM_MPORT_573_en = reset;
  assign RAM_MPORT_574_data = 32'h0;
  assign RAM_MPORT_574_addr = 10'h23e;
  assign RAM_MPORT_574_mask = 1'h1;
  assign RAM_MPORT_574_en = reset;
  assign RAM_MPORT_575_data = 32'h0;
  assign RAM_MPORT_575_addr = 10'h23f;
  assign RAM_MPORT_575_mask = 1'h1;
  assign RAM_MPORT_575_en = reset;
  assign RAM_MPORT_576_data = 32'h0;
  assign RAM_MPORT_576_addr = 10'h240;
  assign RAM_MPORT_576_mask = 1'h1;
  assign RAM_MPORT_576_en = reset;
  assign RAM_MPORT_577_data = 32'h0;
  assign RAM_MPORT_577_addr = 10'h241;
  assign RAM_MPORT_577_mask = 1'h1;
  assign RAM_MPORT_577_en = reset;
  assign RAM_MPORT_578_data = 32'h0;
  assign RAM_MPORT_578_addr = 10'h242;
  assign RAM_MPORT_578_mask = 1'h1;
  assign RAM_MPORT_578_en = reset;
  assign RAM_MPORT_579_data = 32'h0;
  assign RAM_MPORT_579_addr = 10'h243;
  assign RAM_MPORT_579_mask = 1'h1;
  assign RAM_MPORT_579_en = reset;
  assign RAM_MPORT_580_data = 32'h0;
  assign RAM_MPORT_580_addr = 10'h244;
  assign RAM_MPORT_580_mask = 1'h1;
  assign RAM_MPORT_580_en = reset;
  assign RAM_MPORT_581_data = 32'h0;
  assign RAM_MPORT_581_addr = 10'h245;
  assign RAM_MPORT_581_mask = 1'h1;
  assign RAM_MPORT_581_en = reset;
  assign RAM_MPORT_582_data = 32'h0;
  assign RAM_MPORT_582_addr = 10'h246;
  assign RAM_MPORT_582_mask = 1'h1;
  assign RAM_MPORT_582_en = reset;
  assign RAM_MPORT_583_data = 32'h0;
  assign RAM_MPORT_583_addr = 10'h247;
  assign RAM_MPORT_583_mask = 1'h1;
  assign RAM_MPORT_583_en = reset;
  assign RAM_MPORT_584_data = 32'h0;
  assign RAM_MPORT_584_addr = 10'h248;
  assign RAM_MPORT_584_mask = 1'h1;
  assign RAM_MPORT_584_en = reset;
  assign RAM_MPORT_585_data = 32'h0;
  assign RAM_MPORT_585_addr = 10'h249;
  assign RAM_MPORT_585_mask = 1'h1;
  assign RAM_MPORT_585_en = reset;
  assign RAM_MPORT_586_data = 32'h0;
  assign RAM_MPORT_586_addr = 10'h24a;
  assign RAM_MPORT_586_mask = 1'h1;
  assign RAM_MPORT_586_en = reset;
  assign RAM_MPORT_587_data = 32'h0;
  assign RAM_MPORT_587_addr = 10'h24b;
  assign RAM_MPORT_587_mask = 1'h1;
  assign RAM_MPORT_587_en = reset;
  assign RAM_MPORT_588_data = 32'h0;
  assign RAM_MPORT_588_addr = 10'h24c;
  assign RAM_MPORT_588_mask = 1'h1;
  assign RAM_MPORT_588_en = reset;
  assign RAM_MPORT_589_data = 32'h0;
  assign RAM_MPORT_589_addr = 10'h24d;
  assign RAM_MPORT_589_mask = 1'h1;
  assign RAM_MPORT_589_en = reset;
  assign RAM_MPORT_590_data = 32'h0;
  assign RAM_MPORT_590_addr = 10'h24e;
  assign RAM_MPORT_590_mask = 1'h1;
  assign RAM_MPORT_590_en = reset;
  assign RAM_MPORT_591_data = 32'h0;
  assign RAM_MPORT_591_addr = 10'h24f;
  assign RAM_MPORT_591_mask = 1'h1;
  assign RAM_MPORT_591_en = reset;
  assign RAM_MPORT_592_data = 32'h0;
  assign RAM_MPORT_592_addr = 10'h250;
  assign RAM_MPORT_592_mask = 1'h1;
  assign RAM_MPORT_592_en = reset;
  assign RAM_MPORT_593_data = 32'h0;
  assign RAM_MPORT_593_addr = 10'h251;
  assign RAM_MPORT_593_mask = 1'h1;
  assign RAM_MPORT_593_en = reset;
  assign RAM_MPORT_594_data = 32'h0;
  assign RAM_MPORT_594_addr = 10'h252;
  assign RAM_MPORT_594_mask = 1'h1;
  assign RAM_MPORT_594_en = reset;
  assign RAM_MPORT_595_data = 32'h0;
  assign RAM_MPORT_595_addr = 10'h253;
  assign RAM_MPORT_595_mask = 1'h1;
  assign RAM_MPORT_595_en = reset;
  assign RAM_MPORT_596_data = 32'h0;
  assign RAM_MPORT_596_addr = 10'h254;
  assign RAM_MPORT_596_mask = 1'h1;
  assign RAM_MPORT_596_en = reset;
  assign RAM_MPORT_597_data = 32'h0;
  assign RAM_MPORT_597_addr = 10'h255;
  assign RAM_MPORT_597_mask = 1'h1;
  assign RAM_MPORT_597_en = reset;
  assign RAM_MPORT_598_data = 32'h0;
  assign RAM_MPORT_598_addr = 10'h256;
  assign RAM_MPORT_598_mask = 1'h1;
  assign RAM_MPORT_598_en = reset;
  assign RAM_MPORT_599_data = 32'h0;
  assign RAM_MPORT_599_addr = 10'h257;
  assign RAM_MPORT_599_mask = 1'h1;
  assign RAM_MPORT_599_en = reset;
  assign RAM_MPORT_600_data = 32'h0;
  assign RAM_MPORT_600_addr = 10'h258;
  assign RAM_MPORT_600_mask = 1'h1;
  assign RAM_MPORT_600_en = reset;
  assign RAM_MPORT_601_data = 32'h0;
  assign RAM_MPORT_601_addr = 10'h259;
  assign RAM_MPORT_601_mask = 1'h1;
  assign RAM_MPORT_601_en = reset;
  assign RAM_MPORT_602_data = 32'h0;
  assign RAM_MPORT_602_addr = 10'h25a;
  assign RAM_MPORT_602_mask = 1'h1;
  assign RAM_MPORT_602_en = reset;
  assign RAM_MPORT_603_data = 32'h0;
  assign RAM_MPORT_603_addr = 10'h25b;
  assign RAM_MPORT_603_mask = 1'h1;
  assign RAM_MPORT_603_en = reset;
  assign RAM_MPORT_604_data = 32'h0;
  assign RAM_MPORT_604_addr = 10'h25c;
  assign RAM_MPORT_604_mask = 1'h1;
  assign RAM_MPORT_604_en = reset;
  assign RAM_MPORT_605_data = 32'h0;
  assign RAM_MPORT_605_addr = 10'h25d;
  assign RAM_MPORT_605_mask = 1'h1;
  assign RAM_MPORT_605_en = reset;
  assign RAM_MPORT_606_data = 32'h0;
  assign RAM_MPORT_606_addr = 10'h25e;
  assign RAM_MPORT_606_mask = 1'h1;
  assign RAM_MPORT_606_en = reset;
  assign RAM_MPORT_607_data = 32'h0;
  assign RAM_MPORT_607_addr = 10'h25f;
  assign RAM_MPORT_607_mask = 1'h1;
  assign RAM_MPORT_607_en = reset;
  assign RAM_MPORT_608_data = 32'h0;
  assign RAM_MPORT_608_addr = 10'h260;
  assign RAM_MPORT_608_mask = 1'h1;
  assign RAM_MPORT_608_en = reset;
  assign RAM_MPORT_609_data = 32'h0;
  assign RAM_MPORT_609_addr = 10'h261;
  assign RAM_MPORT_609_mask = 1'h1;
  assign RAM_MPORT_609_en = reset;
  assign RAM_MPORT_610_data = 32'h0;
  assign RAM_MPORT_610_addr = 10'h262;
  assign RAM_MPORT_610_mask = 1'h1;
  assign RAM_MPORT_610_en = reset;
  assign RAM_MPORT_611_data = 32'h0;
  assign RAM_MPORT_611_addr = 10'h263;
  assign RAM_MPORT_611_mask = 1'h1;
  assign RAM_MPORT_611_en = reset;
  assign RAM_MPORT_612_data = 32'h0;
  assign RAM_MPORT_612_addr = 10'h264;
  assign RAM_MPORT_612_mask = 1'h1;
  assign RAM_MPORT_612_en = reset;
  assign RAM_MPORT_613_data = 32'h0;
  assign RAM_MPORT_613_addr = 10'h265;
  assign RAM_MPORT_613_mask = 1'h1;
  assign RAM_MPORT_613_en = reset;
  assign RAM_MPORT_614_data = 32'h0;
  assign RAM_MPORT_614_addr = 10'h266;
  assign RAM_MPORT_614_mask = 1'h1;
  assign RAM_MPORT_614_en = reset;
  assign RAM_MPORT_615_data = 32'h0;
  assign RAM_MPORT_615_addr = 10'h267;
  assign RAM_MPORT_615_mask = 1'h1;
  assign RAM_MPORT_615_en = reset;
  assign RAM_MPORT_616_data = 32'h0;
  assign RAM_MPORT_616_addr = 10'h268;
  assign RAM_MPORT_616_mask = 1'h1;
  assign RAM_MPORT_616_en = reset;
  assign RAM_MPORT_617_data = 32'h0;
  assign RAM_MPORT_617_addr = 10'h269;
  assign RAM_MPORT_617_mask = 1'h1;
  assign RAM_MPORT_617_en = reset;
  assign RAM_MPORT_618_data = 32'h0;
  assign RAM_MPORT_618_addr = 10'h26a;
  assign RAM_MPORT_618_mask = 1'h1;
  assign RAM_MPORT_618_en = reset;
  assign RAM_MPORT_619_data = 32'h0;
  assign RAM_MPORT_619_addr = 10'h26b;
  assign RAM_MPORT_619_mask = 1'h1;
  assign RAM_MPORT_619_en = reset;
  assign RAM_MPORT_620_data = 32'h0;
  assign RAM_MPORT_620_addr = 10'h26c;
  assign RAM_MPORT_620_mask = 1'h1;
  assign RAM_MPORT_620_en = reset;
  assign RAM_MPORT_621_data = 32'h0;
  assign RAM_MPORT_621_addr = 10'h26d;
  assign RAM_MPORT_621_mask = 1'h1;
  assign RAM_MPORT_621_en = reset;
  assign RAM_MPORT_622_data = 32'h0;
  assign RAM_MPORT_622_addr = 10'h26e;
  assign RAM_MPORT_622_mask = 1'h1;
  assign RAM_MPORT_622_en = reset;
  assign RAM_MPORT_623_data = 32'h0;
  assign RAM_MPORT_623_addr = 10'h26f;
  assign RAM_MPORT_623_mask = 1'h1;
  assign RAM_MPORT_623_en = reset;
  assign RAM_MPORT_624_data = 32'h0;
  assign RAM_MPORT_624_addr = 10'h270;
  assign RAM_MPORT_624_mask = 1'h1;
  assign RAM_MPORT_624_en = reset;
  assign RAM_MPORT_625_data = 32'h0;
  assign RAM_MPORT_625_addr = 10'h271;
  assign RAM_MPORT_625_mask = 1'h1;
  assign RAM_MPORT_625_en = reset;
  assign RAM_MPORT_626_data = 32'h0;
  assign RAM_MPORT_626_addr = 10'h272;
  assign RAM_MPORT_626_mask = 1'h1;
  assign RAM_MPORT_626_en = reset;
  assign RAM_MPORT_627_data = 32'h0;
  assign RAM_MPORT_627_addr = 10'h273;
  assign RAM_MPORT_627_mask = 1'h1;
  assign RAM_MPORT_627_en = reset;
  assign RAM_MPORT_628_data = 32'h0;
  assign RAM_MPORT_628_addr = 10'h274;
  assign RAM_MPORT_628_mask = 1'h1;
  assign RAM_MPORT_628_en = reset;
  assign RAM_MPORT_629_data = 32'h0;
  assign RAM_MPORT_629_addr = 10'h275;
  assign RAM_MPORT_629_mask = 1'h1;
  assign RAM_MPORT_629_en = reset;
  assign RAM_MPORT_630_data = 32'h0;
  assign RAM_MPORT_630_addr = 10'h276;
  assign RAM_MPORT_630_mask = 1'h1;
  assign RAM_MPORT_630_en = reset;
  assign RAM_MPORT_631_data = 32'h0;
  assign RAM_MPORT_631_addr = 10'h277;
  assign RAM_MPORT_631_mask = 1'h1;
  assign RAM_MPORT_631_en = reset;
  assign RAM_MPORT_632_data = 32'h0;
  assign RAM_MPORT_632_addr = 10'h278;
  assign RAM_MPORT_632_mask = 1'h1;
  assign RAM_MPORT_632_en = reset;
  assign RAM_MPORT_633_data = 32'h0;
  assign RAM_MPORT_633_addr = 10'h279;
  assign RAM_MPORT_633_mask = 1'h1;
  assign RAM_MPORT_633_en = reset;
  assign RAM_MPORT_634_data = 32'h0;
  assign RAM_MPORT_634_addr = 10'h27a;
  assign RAM_MPORT_634_mask = 1'h1;
  assign RAM_MPORT_634_en = reset;
  assign RAM_MPORT_635_data = 32'h0;
  assign RAM_MPORT_635_addr = 10'h27b;
  assign RAM_MPORT_635_mask = 1'h1;
  assign RAM_MPORT_635_en = reset;
  assign RAM_MPORT_636_data = 32'h0;
  assign RAM_MPORT_636_addr = 10'h27c;
  assign RAM_MPORT_636_mask = 1'h1;
  assign RAM_MPORT_636_en = reset;
  assign RAM_MPORT_637_data = 32'h0;
  assign RAM_MPORT_637_addr = 10'h27d;
  assign RAM_MPORT_637_mask = 1'h1;
  assign RAM_MPORT_637_en = reset;
  assign RAM_MPORT_638_data = 32'h0;
  assign RAM_MPORT_638_addr = 10'h27e;
  assign RAM_MPORT_638_mask = 1'h1;
  assign RAM_MPORT_638_en = reset;
  assign RAM_MPORT_639_data = 32'h0;
  assign RAM_MPORT_639_addr = 10'h27f;
  assign RAM_MPORT_639_mask = 1'h1;
  assign RAM_MPORT_639_en = reset;
  assign RAM_MPORT_640_data = 32'h0;
  assign RAM_MPORT_640_addr = 10'h280;
  assign RAM_MPORT_640_mask = 1'h1;
  assign RAM_MPORT_640_en = reset;
  assign RAM_MPORT_641_data = 32'h0;
  assign RAM_MPORT_641_addr = 10'h281;
  assign RAM_MPORT_641_mask = 1'h1;
  assign RAM_MPORT_641_en = reset;
  assign RAM_MPORT_642_data = 32'h0;
  assign RAM_MPORT_642_addr = 10'h282;
  assign RAM_MPORT_642_mask = 1'h1;
  assign RAM_MPORT_642_en = reset;
  assign RAM_MPORT_643_data = 32'h0;
  assign RAM_MPORT_643_addr = 10'h283;
  assign RAM_MPORT_643_mask = 1'h1;
  assign RAM_MPORT_643_en = reset;
  assign RAM_MPORT_644_data = 32'h0;
  assign RAM_MPORT_644_addr = 10'h284;
  assign RAM_MPORT_644_mask = 1'h1;
  assign RAM_MPORT_644_en = reset;
  assign RAM_MPORT_645_data = 32'h0;
  assign RAM_MPORT_645_addr = 10'h285;
  assign RAM_MPORT_645_mask = 1'h1;
  assign RAM_MPORT_645_en = reset;
  assign RAM_MPORT_646_data = 32'h0;
  assign RAM_MPORT_646_addr = 10'h286;
  assign RAM_MPORT_646_mask = 1'h1;
  assign RAM_MPORT_646_en = reset;
  assign RAM_MPORT_647_data = 32'h0;
  assign RAM_MPORT_647_addr = 10'h287;
  assign RAM_MPORT_647_mask = 1'h1;
  assign RAM_MPORT_647_en = reset;
  assign RAM_MPORT_648_data = 32'h0;
  assign RAM_MPORT_648_addr = 10'h288;
  assign RAM_MPORT_648_mask = 1'h1;
  assign RAM_MPORT_648_en = reset;
  assign RAM_MPORT_649_data = 32'h0;
  assign RAM_MPORT_649_addr = 10'h289;
  assign RAM_MPORT_649_mask = 1'h1;
  assign RAM_MPORT_649_en = reset;
  assign RAM_MPORT_650_data = 32'h0;
  assign RAM_MPORT_650_addr = 10'h28a;
  assign RAM_MPORT_650_mask = 1'h1;
  assign RAM_MPORT_650_en = reset;
  assign RAM_MPORT_651_data = 32'h0;
  assign RAM_MPORT_651_addr = 10'h28b;
  assign RAM_MPORT_651_mask = 1'h1;
  assign RAM_MPORT_651_en = reset;
  assign RAM_MPORT_652_data = 32'h0;
  assign RAM_MPORT_652_addr = 10'h28c;
  assign RAM_MPORT_652_mask = 1'h1;
  assign RAM_MPORT_652_en = reset;
  assign RAM_MPORT_653_data = 32'h0;
  assign RAM_MPORT_653_addr = 10'h28d;
  assign RAM_MPORT_653_mask = 1'h1;
  assign RAM_MPORT_653_en = reset;
  assign RAM_MPORT_654_data = 32'h0;
  assign RAM_MPORT_654_addr = 10'h28e;
  assign RAM_MPORT_654_mask = 1'h1;
  assign RAM_MPORT_654_en = reset;
  assign RAM_MPORT_655_data = 32'h0;
  assign RAM_MPORT_655_addr = 10'h28f;
  assign RAM_MPORT_655_mask = 1'h1;
  assign RAM_MPORT_655_en = reset;
  assign RAM_MPORT_656_data = 32'h0;
  assign RAM_MPORT_656_addr = 10'h290;
  assign RAM_MPORT_656_mask = 1'h1;
  assign RAM_MPORT_656_en = reset;
  assign RAM_MPORT_657_data = 32'h0;
  assign RAM_MPORT_657_addr = 10'h291;
  assign RAM_MPORT_657_mask = 1'h1;
  assign RAM_MPORT_657_en = reset;
  assign RAM_MPORT_658_data = 32'h0;
  assign RAM_MPORT_658_addr = 10'h292;
  assign RAM_MPORT_658_mask = 1'h1;
  assign RAM_MPORT_658_en = reset;
  assign RAM_MPORT_659_data = 32'h0;
  assign RAM_MPORT_659_addr = 10'h293;
  assign RAM_MPORT_659_mask = 1'h1;
  assign RAM_MPORT_659_en = reset;
  assign RAM_MPORT_660_data = 32'h0;
  assign RAM_MPORT_660_addr = 10'h294;
  assign RAM_MPORT_660_mask = 1'h1;
  assign RAM_MPORT_660_en = reset;
  assign RAM_MPORT_661_data = 32'h0;
  assign RAM_MPORT_661_addr = 10'h295;
  assign RAM_MPORT_661_mask = 1'h1;
  assign RAM_MPORT_661_en = reset;
  assign RAM_MPORT_662_data = 32'h0;
  assign RAM_MPORT_662_addr = 10'h296;
  assign RAM_MPORT_662_mask = 1'h1;
  assign RAM_MPORT_662_en = reset;
  assign RAM_MPORT_663_data = 32'h0;
  assign RAM_MPORT_663_addr = 10'h297;
  assign RAM_MPORT_663_mask = 1'h1;
  assign RAM_MPORT_663_en = reset;
  assign RAM_MPORT_664_data = 32'h0;
  assign RAM_MPORT_664_addr = 10'h298;
  assign RAM_MPORT_664_mask = 1'h1;
  assign RAM_MPORT_664_en = reset;
  assign RAM_MPORT_665_data = 32'h0;
  assign RAM_MPORT_665_addr = 10'h299;
  assign RAM_MPORT_665_mask = 1'h1;
  assign RAM_MPORT_665_en = reset;
  assign RAM_MPORT_666_data = 32'h0;
  assign RAM_MPORT_666_addr = 10'h29a;
  assign RAM_MPORT_666_mask = 1'h1;
  assign RAM_MPORT_666_en = reset;
  assign RAM_MPORT_667_data = 32'h0;
  assign RAM_MPORT_667_addr = 10'h29b;
  assign RAM_MPORT_667_mask = 1'h1;
  assign RAM_MPORT_667_en = reset;
  assign RAM_MPORT_668_data = 32'h0;
  assign RAM_MPORT_668_addr = 10'h29c;
  assign RAM_MPORT_668_mask = 1'h1;
  assign RAM_MPORT_668_en = reset;
  assign RAM_MPORT_669_data = 32'h0;
  assign RAM_MPORT_669_addr = 10'h29d;
  assign RAM_MPORT_669_mask = 1'h1;
  assign RAM_MPORT_669_en = reset;
  assign RAM_MPORT_670_data = 32'h0;
  assign RAM_MPORT_670_addr = 10'h29e;
  assign RAM_MPORT_670_mask = 1'h1;
  assign RAM_MPORT_670_en = reset;
  assign RAM_MPORT_671_data = 32'h0;
  assign RAM_MPORT_671_addr = 10'h29f;
  assign RAM_MPORT_671_mask = 1'h1;
  assign RAM_MPORT_671_en = reset;
  assign RAM_MPORT_672_data = 32'h0;
  assign RAM_MPORT_672_addr = 10'h2a0;
  assign RAM_MPORT_672_mask = 1'h1;
  assign RAM_MPORT_672_en = reset;
  assign RAM_MPORT_673_data = 32'h0;
  assign RAM_MPORT_673_addr = 10'h2a1;
  assign RAM_MPORT_673_mask = 1'h1;
  assign RAM_MPORT_673_en = reset;
  assign RAM_MPORT_674_data = 32'h0;
  assign RAM_MPORT_674_addr = 10'h2a2;
  assign RAM_MPORT_674_mask = 1'h1;
  assign RAM_MPORT_674_en = reset;
  assign RAM_MPORT_675_data = 32'h0;
  assign RAM_MPORT_675_addr = 10'h2a3;
  assign RAM_MPORT_675_mask = 1'h1;
  assign RAM_MPORT_675_en = reset;
  assign RAM_MPORT_676_data = 32'h0;
  assign RAM_MPORT_676_addr = 10'h2a4;
  assign RAM_MPORT_676_mask = 1'h1;
  assign RAM_MPORT_676_en = reset;
  assign RAM_MPORT_677_data = 32'h0;
  assign RAM_MPORT_677_addr = 10'h2a5;
  assign RAM_MPORT_677_mask = 1'h1;
  assign RAM_MPORT_677_en = reset;
  assign RAM_MPORT_678_data = 32'h0;
  assign RAM_MPORT_678_addr = 10'h2a6;
  assign RAM_MPORT_678_mask = 1'h1;
  assign RAM_MPORT_678_en = reset;
  assign RAM_MPORT_679_data = 32'h0;
  assign RAM_MPORT_679_addr = 10'h2a7;
  assign RAM_MPORT_679_mask = 1'h1;
  assign RAM_MPORT_679_en = reset;
  assign RAM_MPORT_680_data = 32'h0;
  assign RAM_MPORT_680_addr = 10'h2a8;
  assign RAM_MPORT_680_mask = 1'h1;
  assign RAM_MPORT_680_en = reset;
  assign RAM_MPORT_681_data = 32'h0;
  assign RAM_MPORT_681_addr = 10'h2a9;
  assign RAM_MPORT_681_mask = 1'h1;
  assign RAM_MPORT_681_en = reset;
  assign RAM_MPORT_682_data = 32'h0;
  assign RAM_MPORT_682_addr = 10'h2aa;
  assign RAM_MPORT_682_mask = 1'h1;
  assign RAM_MPORT_682_en = reset;
  assign RAM_MPORT_683_data = 32'h0;
  assign RAM_MPORT_683_addr = 10'h2ab;
  assign RAM_MPORT_683_mask = 1'h1;
  assign RAM_MPORT_683_en = reset;
  assign RAM_MPORT_684_data = 32'h0;
  assign RAM_MPORT_684_addr = 10'h2ac;
  assign RAM_MPORT_684_mask = 1'h1;
  assign RAM_MPORT_684_en = reset;
  assign RAM_MPORT_685_data = 32'h0;
  assign RAM_MPORT_685_addr = 10'h2ad;
  assign RAM_MPORT_685_mask = 1'h1;
  assign RAM_MPORT_685_en = reset;
  assign RAM_MPORT_686_data = 32'h0;
  assign RAM_MPORT_686_addr = 10'h2ae;
  assign RAM_MPORT_686_mask = 1'h1;
  assign RAM_MPORT_686_en = reset;
  assign RAM_MPORT_687_data = 32'h0;
  assign RAM_MPORT_687_addr = 10'h2af;
  assign RAM_MPORT_687_mask = 1'h1;
  assign RAM_MPORT_687_en = reset;
  assign RAM_MPORT_688_data = 32'h0;
  assign RAM_MPORT_688_addr = 10'h2b0;
  assign RAM_MPORT_688_mask = 1'h1;
  assign RAM_MPORT_688_en = reset;
  assign RAM_MPORT_689_data = 32'h0;
  assign RAM_MPORT_689_addr = 10'h2b1;
  assign RAM_MPORT_689_mask = 1'h1;
  assign RAM_MPORT_689_en = reset;
  assign RAM_MPORT_690_data = 32'h0;
  assign RAM_MPORT_690_addr = 10'h2b2;
  assign RAM_MPORT_690_mask = 1'h1;
  assign RAM_MPORT_690_en = reset;
  assign RAM_MPORT_691_data = 32'h0;
  assign RAM_MPORT_691_addr = 10'h2b3;
  assign RAM_MPORT_691_mask = 1'h1;
  assign RAM_MPORT_691_en = reset;
  assign RAM_MPORT_692_data = 32'h0;
  assign RAM_MPORT_692_addr = 10'h2b4;
  assign RAM_MPORT_692_mask = 1'h1;
  assign RAM_MPORT_692_en = reset;
  assign RAM_MPORT_693_data = 32'h0;
  assign RAM_MPORT_693_addr = 10'h2b5;
  assign RAM_MPORT_693_mask = 1'h1;
  assign RAM_MPORT_693_en = reset;
  assign RAM_MPORT_694_data = 32'h0;
  assign RAM_MPORT_694_addr = 10'h2b6;
  assign RAM_MPORT_694_mask = 1'h1;
  assign RAM_MPORT_694_en = reset;
  assign RAM_MPORT_695_data = 32'h0;
  assign RAM_MPORT_695_addr = 10'h2b7;
  assign RAM_MPORT_695_mask = 1'h1;
  assign RAM_MPORT_695_en = reset;
  assign RAM_MPORT_696_data = 32'h0;
  assign RAM_MPORT_696_addr = 10'h2b8;
  assign RAM_MPORT_696_mask = 1'h1;
  assign RAM_MPORT_696_en = reset;
  assign RAM_MPORT_697_data = 32'h0;
  assign RAM_MPORT_697_addr = 10'h2b9;
  assign RAM_MPORT_697_mask = 1'h1;
  assign RAM_MPORT_697_en = reset;
  assign RAM_MPORT_698_data = 32'h0;
  assign RAM_MPORT_698_addr = 10'h2ba;
  assign RAM_MPORT_698_mask = 1'h1;
  assign RAM_MPORT_698_en = reset;
  assign RAM_MPORT_699_data = 32'h0;
  assign RAM_MPORT_699_addr = 10'h2bb;
  assign RAM_MPORT_699_mask = 1'h1;
  assign RAM_MPORT_699_en = reset;
  assign RAM_MPORT_700_data = 32'h0;
  assign RAM_MPORT_700_addr = 10'h2bc;
  assign RAM_MPORT_700_mask = 1'h1;
  assign RAM_MPORT_700_en = reset;
  assign RAM_MPORT_701_data = 32'h0;
  assign RAM_MPORT_701_addr = 10'h2bd;
  assign RAM_MPORT_701_mask = 1'h1;
  assign RAM_MPORT_701_en = reset;
  assign RAM_MPORT_702_data = 32'h0;
  assign RAM_MPORT_702_addr = 10'h2be;
  assign RAM_MPORT_702_mask = 1'h1;
  assign RAM_MPORT_702_en = reset;
  assign RAM_MPORT_703_data = 32'h0;
  assign RAM_MPORT_703_addr = 10'h2bf;
  assign RAM_MPORT_703_mask = 1'h1;
  assign RAM_MPORT_703_en = reset;
  assign RAM_MPORT_704_data = 32'h0;
  assign RAM_MPORT_704_addr = 10'h2c0;
  assign RAM_MPORT_704_mask = 1'h1;
  assign RAM_MPORT_704_en = reset;
  assign RAM_MPORT_705_data = 32'h0;
  assign RAM_MPORT_705_addr = 10'h2c1;
  assign RAM_MPORT_705_mask = 1'h1;
  assign RAM_MPORT_705_en = reset;
  assign RAM_MPORT_706_data = 32'h0;
  assign RAM_MPORT_706_addr = 10'h2c2;
  assign RAM_MPORT_706_mask = 1'h1;
  assign RAM_MPORT_706_en = reset;
  assign RAM_MPORT_707_data = 32'h0;
  assign RAM_MPORT_707_addr = 10'h2c3;
  assign RAM_MPORT_707_mask = 1'h1;
  assign RAM_MPORT_707_en = reset;
  assign RAM_MPORT_708_data = 32'h0;
  assign RAM_MPORT_708_addr = 10'h2c4;
  assign RAM_MPORT_708_mask = 1'h1;
  assign RAM_MPORT_708_en = reset;
  assign RAM_MPORT_709_data = 32'h0;
  assign RAM_MPORT_709_addr = 10'h2c5;
  assign RAM_MPORT_709_mask = 1'h1;
  assign RAM_MPORT_709_en = reset;
  assign RAM_MPORT_710_data = 32'h0;
  assign RAM_MPORT_710_addr = 10'h2c6;
  assign RAM_MPORT_710_mask = 1'h1;
  assign RAM_MPORT_710_en = reset;
  assign RAM_MPORT_711_data = 32'h0;
  assign RAM_MPORT_711_addr = 10'h2c7;
  assign RAM_MPORT_711_mask = 1'h1;
  assign RAM_MPORT_711_en = reset;
  assign RAM_MPORT_712_data = 32'h0;
  assign RAM_MPORT_712_addr = 10'h2c8;
  assign RAM_MPORT_712_mask = 1'h1;
  assign RAM_MPORT_712_en = reset;
  assign RAM_MPORT_713_data = 32'h0;
  assign RAM_MPORT_713_addr = 10'h2c9;
  assign RAM_MPORT_713_mask = 1'h1;
  assign RAM_MPORT_713_en = reset;
  assign RAM_MPORT_714_data = 32'h0;
  assign RAM_MPORT_714_addr = 10'h2ca;
  assign RAM_MPORT_714_mask = 1'h1;
  assign RAM_MPORT_714_en = reset;
  assign RAM_MPORT_715_data = 32'h0;
  assign RAM_MPORT_715_addr = 10'h2cb;
  assign RAM_MPORT_715_mask = 1'h1;
  assign RAM_MPORT_715_en = reset;
  assign RAM_MPORT_716_data = 32'h0;
  assign RAM_MPORT_716_addr = 10'h2cc;
  assign RAM_MPORT_716_mask = 1'h1;
  assign RAM_MPORT_716_en = reset;
  assign RAM_MPORT_717_data = 32'h0;
  assign RAM_MPORT_717_addr = 10'h2cd;
  assign RAM_MPORT_717_mask = 1'h1;
  assign RAM_MPORT_717_en = reset;
  assign RAM_MPORT_718_data = 32'h0;
  assign RAM_MPORT_718_addr = 10'h2ce;
  assign RAM_MPORT_718_mask = 1'h1;
  assign RAM_MPORT_718_en = reset;
  assign RAM_MPORT_719_data = 32'h0;
  assign RAM_MPORT_719_addr = 10'h2cf;
  assign RAM_MPORT_719_mask = 1'h1;
  assign RAM_MPORT_719_en = reset;
  assign RAM_MPORT_720_data = 32'h0;
  assign RAM_MPORT_720_addr = 10'h2d0;
  assign RAM_MPORT_720_mask = 1'h1;
  assign RAM_MPORT_720_en = reset;
  assign RAM_MPORT_721_data = 32'h0;
  assign RAM_MPORT_721_addr = 10'h2d1;
  assign RAM_MPORT_721_mask = 1'h1;
  assign RAM_MPORT_721_en = reset;
  assign RAM_MPORT_722_data = 32'h0;
  assign RAM_MPORT_722_addr = 10'h2d2;
  assign RAM_MPORT_722_mask = 1'h1;
  assign RAM_MPORT_722_en = reset;
  assign RAM_MPORT_723_data = 32'h0;
  assign RAM_MPORT_723_addr = 10'h2d3;
  assign RAM_MPORT_723_mask = 1'h1;
  assign RAM_MPORT_723_en = reset;
  assign RAM_MPORT_724_data = 32'h0;
  assign RAM_MPORT_724_addr = 10'h2d4;
  assign RAM_MPORT_724_mask = 1'h1;
  assign RAM_MPORT_724_en = reset;
  assign RAM_MPORT_725_data = 32'h0;
  assign RAM_MPORT_725_addr = 10'h2d5;
  assign RAM_MPORT_725_mask = 1'h1;
  assign RAM_MPORT_725_en = reset;
  assign RAM_MPORT_726_data = 32'h0;
  assign RAM_MPORT_726_addr = 10'h2d6;
  assign RAM_MPORT_726_mask = 1'h1;
  assign RAM_MPORT_726_en = reset;
  assign RAM_MPORT_727_data = 32'h0;
  assign RAM_MPORT_727_addr = 10'h2d7;
  assign RAM_MPORT_727_mask = 1'h1;
  assign RAM_MPORT_727_en = reset;
  assign RAM_MPORT_728_data = 32'h0;
  assign RAM_MPORT_728_addr = 10'h2d8;
  assign RAM_MPORT_728_mask = 1'h1;
  assign RAM_MPORT_728_en = reset;
  assign RAM_MPORT_729_data = 32'h0;
  assign RAM_MPORT_729_addr = 10'h2d9;
  assign RAM_MPORT_729_mask = 1'h1;
  assign RAM_MPORT_729_en = reset;
  assign RAM_MPORT_730_data = 32'h0;
  assign RAM_MPORT_730_addr = 10'h2da;
  assign RAM_MPORT_730_mask = 1'h1;
  assign RAM_MPORT_730_en = reset;
  assign RAM_MPORT_731_data = 32'h0;
  assign RAM_MPORT_731_addr = 10'h2db;
  assign RAM_MPORT_731_mask = 1'h1;
  assign RAM_MPORT_731_en = reset;
  assign RAM_MPORT_732_data = 32'h0;
  assign RAM_MPORT_732_addr = 10'h2dc;
  assign RAM_MPORT_732_mask = 1'h1;
  assign RAM_MPORT_732_en = reset;
  assign RAM_MPORT_733_data = 32'h0;
  assign RAM_MPORT_733_addr = 10'h2dd;
  assign RAM_MPORT_733_mask = 1'h1;
  assign RAM_MPORT_733_en = reset;
  assign RAM_MPORT_734_data = 32'h0;
  assign RAM_MPORT_734_addr = 10'h2de;
  assign RAM_MPORT_734_mask = 1'h1;
  assign RAM_MPORT_734_en = reset;
  assign RAM_MPORT_735_data = 32'h0;
  assign RAM_MPORT_735_addr = 10'h2df;
  assign RAM_MPORT_735_mask = 1'h1;
  assign RAM_MPORT_735_en = reset;
  assign RAM_MPORT_736_data = 32'h0;
  assign RAM_MPORT_736_addr = 10'h2e0;
  assign RAM_MPORT_736_mask = 1'h1;
  assign RAM_MPORT_736_en = reset;
  assign RAM_MPORT_737_data = 32'h0;
  assign RAM_MPORT_737_addr = 10'h2e1;
  assign RAM_MPORT_737_mask = 1'h1;
  assign RAM_MPORT_737_en = reset;
  assign RAM_MPORT_738_data = 32'h0;
  assign RAM_MPORT_738_addr = 10'h2e2;
  assign RAM_MPORT_738_mask = 1'h1;
  assign RAM_MPORT_738_en = reset;
  assign RAM_MPORT_739_data = 32'h0;
  assign RAM_MPORT_739_addr = 10'h2e3;
  assign RAM_MPORT_739_mask = 1'h1;
  assign RAM_MPORT_739_en = reset;
  assign RAM_MPORT_740_data = 32'h0;
  assign RAM_MPORT_740_addr = 10'h2e4;
  assign RAM_MPORT_740_mask = 1'h1;
  assign RAM_MPORT_740_en = reset;
  assign RAM_MPORT_741_data = 32'h0;
  assign RAM_MPORT_741_addr = 10'h2e5;
  assign RAM_MPORT_741_mask = 1'h1;
  assign RAM_MPORT_741_en = reset;
  assign RAM_MPORT_742_data = 32'h0;
  assign RAM_MPORT_742_addr = 10'h2e6;
  assign RAM_MPORT_742_mask = 1'h1;
  assign RAM_MPORT_742_en = reset;
  assign RAM_MPORT_743_data = 32'h0;
  assign RAM_MPORT_743_addr = 10'h2e7;
  assign RAM_MPORT_743_mask = 1'h1;
  assign RAM_MPORT_743_en = reset;
  assign RAM_MPORT_744_data = 32'h0;
  assign RAM_MPORT_744_addr = 10'h2e8;
  assign RAM_MPORT_744_mask = 1'h1;
  assign RAM_MPORT_744_en = reset;
  assign RAM_MPORT_745_data = 32'h0;
  assign RAM_MPORT_745_addr = 10'h2e9;
  assign RAM_MPORT_745_mask = 1'h1;
  assign RAM_MPORT_745_en = reset;
  assign RAM_MPORT_746_data = 32'h0;
  assign RAM_MPORT_746_addr = 10'h2ea;
  assign RAM_MPORT_746_mask = 1'h1;
  assign RAM_MPORT_746_en = reset;
  assign RAM_MPORT_747_data = 32'h0;
  assign RAM_MPORT_747_addr = 10'h2eb;
  assign RAM_MPORT_747_mask = 1'h1;
  assign RAM_MPORT_747_en = reset;
  assign RAM_MPORT_748_data = 32'h0;
  assign RAM_MPORT_748_addr = 10'h2ec;
  assign RAM_MPORT_748_mask = 1'h1;
  assign RAM_MPORT_748_en = reset;
  assign RAM_MPORT_749_data = 32'h0;
  assign RAM_MPORT_749_addr = 10'h2ed;
  assign RAM_MPORT_749_mask = 1'h1;
  assign RAM_MPORT_749_en = reset;
  assign RAM_MPORT_750_data = 32'h0;
  assign RAM_MPORT_750_addr = 10'h2ee;
  assign RAM_MPORT_750_mask = 1'h1;
  assign RAM_MPORT_750_en = reset;
  assign RAM_MPORT_751_data = 32'h0;
  assign RAM_MPORT_751_addr = 10'h2ef;
  assign RAM_MPORT_751_mask = 1'h1;
  assign RAM_MPORT_751_en = reset;
  assign RAM_MPORT_752_data = 32'h0;
  assign RAM_MPORT_752_addr = 10'h2f0;
  assign RAM_MPORT_752_mask = 1'h1;
  assign RAM_MPORT_752_en = reset;
  assign RAM_MPORT_753_data = 32'h0;
  assign RAM_MPORT_753_addr = 10'h2f1;
  assign RAM_MPORT_753_mask = 1'h1;
  assign RAM_MPORT_753_en = reset;
  assign RAM_MPORT_754_data = 32'h0;
  assign RAM_MPORT_754_addr = 10'h2f2;
  assign RAM_MPORT_754_mask = 1'h1;
  assign RAM_MPORT_754_en = reset;
  assign RAM_MPORT_755_data = 32'h0;
  assign RAM_MPORT_755_addr = 10'h2f3;
  assign RAM_MPORT_755_mask = 1'h1;
  assign RAM_MPORT_755_en = reset;
  assign RAM_MPORT_756_data = 32'h0;
  assign RAM_MPORT_756_addr = 10'h2f4;
  assign RAM_MPORT_756_mask = 1'h1;
  assign RAM_MPORT_756_en = reset;
  assign RAM_MPORT_757_data = 32'h0;
  assign RAM_MPORT_757_addr = 10'h2f5;
  assign RAM_MPORT_757_mask = 1'h1;
  assign RAM_MPORT_757_en = reset;
  assign RAM_MPORT_758_data = 32'h0;
  assign RAM_MPORT_758_addr = 10'h2f6;
  assign RAM_MPORT_758_mask = 1'h1;
  assign RAM_MPORT_758_en = reset;
  assign RAM_MPORT_759_data = 32'h0;
  assign RAM_MPORT_759_addr = 10'h2f7;
  assign RAM_MPORT_759_mask = 1'h1;
  assign RAM_MPORT_759_en = reset;
  assign RAM_MPORT_760_data = 32'h0;
  assign RAM_MPORT_760_addr = 10'h2f8;
  assign RAM_MPORT_760_mask = 1'h1;
  assign RAM_MPORT_760_en = reset;
  assign RAM_MPORT_761_data = 32'h0;
  assign RAM_MPORT_761_addr = 10'h2f9;
  assign RAM_MPORT_761_mask = 1'h1;
  assign RAM_MPORT_761_en = reset;
  assign RAM_MPORT_762_data = 32'h0;
  assign RAM_MPORT_762_addr = 10'h2fa;
  assign RAM_MPORT_762_mask = 1'h1;
  assign RAM_MPORT_762_en = reset;
  assign RAM_MPORT_763_data = 32'h0;
  assign RAM_MPORT_763_addr = 10'h2fb;
  assign RAM_MPORT_763_mask = 1'h1;
  assign RAM_MPORT_763_en = reset;
  assign RAM_MPORT_764_data = 32'h0;
  assign RAM_MPORT_764_addr = 10'h2fc;
  assign RAM_MPORT_764_mask = 1'h1;
  assign RAM_MPORT_764_en = reset;
  assign RAM_MPORT_765_data = 32'h0;
  assign RAM_MPORT_765_addr = 10'h2fd;
  assign RAM_MPORT_765_mask = 1'h1;
  assign RAM_MPORT_765_en = reset;
  assign RAM_MPORT_766_data = 32'h0;
  assign RAM_MPORT_766_addr = 10'h2fe;
  assign RAM_MPORT_766_mask = 1'h1;
  assign RAM_MPORT_766_en = reset;
  assign RAM_MPORT_767_data = 32'h0;
  assign RAM_MPORT_767_addr = 10'h2ff;
  assign RAM_MPORT_767_mask = 1'h1;
  assign RAM_MPORT_767_en = reset;
  assign RAM_MPORT_768_data = 32'h0;
  assign RAM_MPORT_768_addr = 10'h300;
  assign RAM_MPORT_768_mask = 1'h1;
  assign RAM_MPORT_768_en = reset;
  assign RAM_MPORT_769_data = 32'h0;
  assign RAM_MPORT_769_addr = 10'h301;
  assign RAM_MPORT_769_mask = 1'h1;
  assign RAM_MPORT_769_en = reset;
  assign RAM_MPORT_770_data = 32'h0;
  assign RAM_MPORT_770_addr = 10'h302;
  assign RAM_MPORT_770_mask = 1'h1;
  assign RAM_MPORT_770_en = reset;
  assign RAM_MPORT_771_data = 32'h0;
  assign RAM_MPORT_771_addr = 10'h303;
  assign RAM_MPORT_771_mask = 1'h1;
  assign RAM_MPORT_771_en = reset;
  assign RAM_MPORT_772_data = 32'h0;
  assign RAM_MPORT_772_addr = 10'h304;
  assign RAM_MPORT_772_mask = 1'h1;
  assign RAM_MPORT_772_en = reset;
  assign RAM_MPORT_773_data = 32'h0;
  assign RAM_MPORT_773_addr = 10'h305;
  assign RAM_MPORT_773_mask = 1'h1;
  assign RAM_MPORT_773_en = reset;
  assign RAM_MPORT_774_data = 32'h0;
  assign RAM_MPORT_774_addr = 10'h306;
  assign RAM_MPORT_774_mask = 1'h1;
  assign RAM_MPORT_774_en = reset;
  assign RAM_MPORT_775_data = 32'h0;
  assign RAM_MPORT_775_addr = 10'h307;
  assign RAM_MPORT_775_mask = 1'h1;
  assign RAM_MPORT_775_en = reset;
  assign RAM_MPORT_776_data = 32'h0;
  assign RAM_MPORT_776_addr = 10'h308;
  assign RAM_MPORT_776_mask = 1'h1;
  assign RAM_MPORT_776_en = reset;
  assign RAM_MPORT_777_data = 32'h0;
  assign RAM_MPORT_777_addr = 10'h309;
  assign RAM_MPORT_777_mask = 1'h1;
  assign RAM_MPORT_777_en = reset;
  assign RAM_MPORT_778_data = 32'h0;
  assign RAM_MPORT_778_addr = 10'h30a;
  assign RAM_MPORT_778_mask = 1'h1;
  assign RAM_MPORT_778_en = reset;
  assign RAM_MPORT_779_data = 32'h0;
  assign RAM_MPORT_779_addr = 10'h30b;
  assign RAM_MPORT_779_mask = 1'h1;
  assign RAM_MPORT_779_en = reset;
  assign RAM_MPORT_780_data = 32'h0;
  assign RAM_MPORT_780_addr = 10'h30c;
  assign RAM_MPORT_780_mask = 1'h1;
  assign RAM_MPORT_780_en = reset;
  assign RAM_MPORT_781_data = 32'h0;
  assign RAM_MPORT_781_addr = 10'h30d;
  assign RAM_MPORT_781_mask = 1'h1;
  assign RAM_MPORT_781_en = reset;
  assign RAM_MPORT_782_data = 32'h0;
  assign RAM_MPORT_782_addr = 10'h30e;
  assign RAM_MPORT_782_mask = 1'h1;
  assign RAM_MPORT_782_en = reset;
  assign RAM_MPORT_783_data = 32'h0;
  assign RAM_MPORT_783_addr = 10'h30f;
  assign RAM_MPORT_783_mask = 1'h1;
  assign RAM_MPORT_783_en = reset;
  assign RAM_MPORT_784_data = 32'h0;
  assign RAM_MPORT_784_addr = 10'h310;
  assign RAM_MPORT_784_mask = 1'h1;
  assign RAM_MPORT_784_en = reset;
  assign RAM_MPORT_785_data = 32'h0;
  assign RAM_MPORT_785_addr = 10'h311;
  assign RAM_MPORT_785_mask = 1'h1;
  assign RAM_MPORT_785_en = reset;
  assign RAM_MPORT_786_data = 32'h0;
  assign RAM_MPORT_786_addr = 10'h312;
  assign RAM_MPORT_786_mask = 1'h1;
  assign RAM_MPORT_786_en = reset;
  assign RAM_MPORT_787_data = 32'h0;
  assign RAM_MPORT_787_addr = 10'h313;
  assign RAM_MPORT_787_mask = 1'h1;
  assign RAM_MPORT_787_en = reset;
  assign RAM_MPORT_788_data = 32'h0;
  assign RAM_MPORT_788_addr = 10'h314;
  assign RAM_MPORT_788_mask = 1'h1;
  assign RAM_MPORT_788_en = reset;
  assign RAM_MPORT_789_data = 32'h0;
  assign RAM_MPORT_789_addr = 10'h315;
  assign RAM_MPORT_789_mask = 1'h1;
  assign RAM_MPORT_789_en = reset;
  assign RAM_MPORT_790_data = 32'h0;
  assign RAM_MPORT_790_addr = 10'h316;
  assign RAM_MPORT_790_mask = 1'h1;
  assign RAM_MPORT_790_en = reset;
  assign RAM_MPORT_791_data = 32'h0;
  assign RAM_MPORT_791_addr = 10'h317;
  assign RAM_MPORT_791_mask = 1'h1;
  assign RAM_MPORT_791_en = reset;
  assign RAM_MPORT_792_data = 32'h0;
  assign RAM_MPORT_792_addr = 10'h318;
  assign RAM_MPORT_792_mask = 1'h1;
  assign RAM_MPORT_792_en = reset;
  assign RAM_MPORT_793_data = 32'h0;
  assign RAM_MPORT_793_addr = 10'h319;
  assign RAM_MPORT_793_mask = 1'h1;
  assign RAM_MPORT_793_en = reset;
  assign RAM_MPORT_794_data = 32'h0;
  assign RAM_MPORT_794_addr = 10'h31a;
  assign RAM_MPORT_794_mask = 1'h1;
  assign RAM_MPORT_794_en = reset;
  assign RAM_MPORT_795_data = 32'h0;
  assign RAM_MPORT_795_addr = 10'h31b;
  assign RAM_MPORT_795_mask = 1'h1;
  assign RAM_MPORT_795_en = reset;
  assign RAM_MPORT_796_data = 32'h0;
  assign RAM_MPORT_796_addr = 10'h31c;
  assign RAM_MPORT_796_mask = 1'h1;
  assign RAM_MPORT_796_en = reset;
  assign RAM_MPORT_797_data = 32'h0;
  assign RAM_MPORT_797_addr = 10'h31d;
  assign RAM_MPORT_797_mask = 1'h1;
  assign RAM_MPORT_797_en = reset;
  assign RAM_MPORT_798_data = 32'h0;
  assign RAM_MPORT_798_addr = 10'h31e;
  assign RAM_MPORT_798_mask = 1'h1;
  assign RAM_MPORT_798_en = reset;
  assign RAM_MPORT_799_data = 32'h0;
  assign RAM_MPORT_799_addr = 10'h31f;
  assign RAM_MPORT_799_mask = 1'h1;
  assign RAM_MPORT_799_en = reset;
  assign RAM_MPORT_800_data = 32'h0;
  assign RAM_MPORT_800_addr = 10'h320;
  assign RAM_MPORT_800_mask = 1'h1;
  assign RAM_MPORT_800_en = reset;
  assign RAM_MPORT_801_data = 32'h0;
  assign RAM_MPORT_801_addr = 10'h321;
  assign RAM_MPORT_801_mask = 1'h1;
  assign RAM_MPORT_801_en = reset;
  assign RAM_MPORT_802_data = 32'h0;
  assign RAM_MPORT_802_addr = 10'h322;
  assign RAM_MPORT_802_mask = 1'h1;
  assign RAM_MPORT_802_en = reset;
  assign RAM_MPORT_803_data = 32'h0;
  assign RAM_MPORT_803_addr = 10'h323;
  assign RAM_MPORT_803_mask = 1'h1;
  assign RAM_MPORT_803_en = reset;
  assign RAM_MPORT_804_data = 32'h0;
  assign RAM_MPORT_804_addr = 10'h324;
  assign RAM_MPORT_804_mask = 1'h1;
  assign RAM_MPORT_804_en = reset;
  assign RAM_MPORT_805_data = 32'h0;
  assign RAM_MPORT_805_addr = 10'h325;
  assign RAM_MPORT_805_mask = 1'h1;
  assign RAM_MPORT_805_en = reset;
  assign RAM_MPORT_806_data = 32'h0;
  assign RAM_MPORT_806_addr = 10'h326;
  assign RAM_MPORT_806_mask = 1'h1;
  assign RAM_MPORT_806_en = reset;
  assign RAM_MPORT_807_data = 32'h0;
  assign RAM_MPORT_807_addr = 10'h327;
  assign RAM_MPORT_807_mask = 1'h1;
  assign RAM_MPORT_807_en = reset;
  assign RAM_MPORT_808_data = 32'h0;
  assign RAM_MPORT_808_addr = 10'h328;
  assign RAM_MPORT_808_mask = 1'h1;
  assign RAM_MPORT_808_en = reset;
  assign RAM_MPORT_809_data = 32'h0;
  assign RAM_MPORT_809_addr = 10'h329;
  assign RAM_MPORT_809_mask = 1'h1;
  assign RAM_MPORT_809_en = reset;
  assign RAM_MPORT_810_data = 32'h0;
  assign RAM_MPORT_810_addr = 10'h32a;
  assign RAM_MPORT_810_mask = 1'h1;
  assign RAM_MPORT_810_en = reset;
  assign RAM_MPORT_811_data = 32'h0;
  assign RAM_MPORT_811_addr = 10'h32b;
  assign RAM_MPORT_811_mask = 1'h1;
  assign RAM_MPORT_811_en = reset;
  assign RAM_MPORT_812_data = 32'h0;
  assign RAM_MPORT_812_addr = 10'h32c;
  assign RAM_MPORT_812_mask = 1'h1;
  assign RAM_MPORT_812_en = reset;
  assign RAM_MPORT_813_data = 32'h0;
  assign RAM_MPORT_813_addr = 10'h32d;
  assign RAM_MPORT_813_mask = 1'h1;
  assign RAM_MPORT_813_en = reset;
  assign RAM_MPORT_814_data = 32'h0;
  assign RAM_MPORT_814_addr = 10'h32e;
  assign RAM_MPORT_814_mask = 1'h1;
  assign RAM_MPORT_814_en = reset;
  assign RAM_MPORT_815_data = 32'h0;
  assign RAM_MPORT_815_addr = 10'h32f;
  assign RAM_MPORT_815_mask = 1'h1;
  assign RAM_MPORT_815_en = reset;
  assign RAM_MPORT_816_data = 32'h0;
  assign RAM_MPORT_816_addr = 10'h330;
  assign RAM_MPORT_816_mask = 1'h1;
  assign RAM_MPORT_816_en = reset;
  assign RAM_MPORT_817_data = 32'h0;
  assign RAM_MPORT_817_addr = 10'h331;
  assign RAM_MPORT_817_mask = 1'h1;
  assign RAM_MPORT_817_en = reset;
  assign RAM_MPORT_818_data = 32'h0;
  assign RAM_MPORT_818_addr = 10'h332;
  assign RAM_MPORT_818_mask = 1'h1;
  assign RAM_MPORT_818_en = reset;
  assign RAM_MPORT_819_data = 32'h0;
  assign RAM_MPORT_819_addr = 10'h333;
  assign RAM_MPORT_819_mask = 1'h1;
  assign RAM_MPORT_819_en = reset;
  assign RAM_MPORT_820_data = 32'h0;
  assign RAM_MPORT_820_addr = 10'h334;
  assign RAM_MPORT_820_mask = 1'h1;
  assign RAM_MPORT_820_en = reset;
  assign RAM_MPORT_821_data = 32'h0;
  assign RAM_MPORT_821_addr = 10'h335;
  assign RAM_MPORT_821_mask = 1'h1;
  assign RAM_MPORT_821_en = reset;
  assign RAM_MPORT_822_data = 32'h0;
  assign RAM_MPORT_822_addr = 10'h336;
  assign RAM_MPORT_822_mask = 1'h1;
  assign RAM_MPORT_822_en = reset;
  assign RAM_MPORT_823_data = 32'h0;
  assign RAM_MPORT_823_addr = 10'h337;
  assign RAM_MPORT_823_mask = 1'h1;
  assign RAM_MPORT_823_en = reset;
  assign RAM_MPORT_824_data = 32'h0;
  assign RAM_MPORT_824_addr = 10'h338;
  assign RAM_MPORT_824_mask = 1'h1;
  assign RAM_MPORT_824_en = reset;
  assign RAM_MPORT_825_data = 32'h0;
  assign RAM_MPORT_825_addr = 10'h339;
  assign RAM_MPORT_825_mask = 1'h1;
  assign RAM_MPORT_825_en = reset;
  assign RAM_MPORT_826_data = 32'h0;
  assign RAM_MPORT_826_addr = 10'h33a;
  assign RAM_MPORT_826_mask = 1'h1;
  assign RAM_MPORT_826_en = reset;
  assign RAM_MPORT_827_data = 32'h0;
  assign RAM_MPORT_827_addr = 10'h33b;
  assign RAM_MPORT_827_mask = 1'h1;
  assign RAM_MPORT_827_en = reset;
  assign RAM_MPORT_828_data = 32'h0;
  assign RAM_MPORT_828_addr = 10'h33c;
  assign RAM_MPORT_828_mask = 1'h1;
  assign RAM_MPORT_828_en = reset;
  assign RAM_MPORT_829_data = 32'h0;
  assign RAM_MPORT_829_addr = 10'h33d;
  assign RAM_MPORT_829_mask = 1'h1;
  assign RAM_MPORT_829_en = reset;
  assign RAM_MPORT_830_data = 32'h0;
  assign RAM_MPORT_830_addr = 10'h33e;
  assign RAM_MPORT_830_mask = 1'h1;
  assign RAM_MPORT_830_en = reset;
  assign RAM_MPORT_831_data = 32'h0;
  assign RAM_MPORT_831_addr = 10'h33f;
  assign RAM_MPORT_831_mask = 1'h1;
  assign RAM_MPORT_831_en = reset;
  assign RAM_MPORT_832_data = 32'h0;
  assign RAM_MPORT_832_addr = 10'h340;
  assign RAM_MPORT_832_mask = 1'h1;
  assign RAM_MPORT_832_en = reset;
  assign RAM_MPORT_833_data = 32'h0;
  assign RAM_MPORT_833_addr = 10'h341;
  assign RAM_MPORT_833_mask = 1'h1;
  assign RAM_MPORT_833_en = reset;
  assign RAM_MPORT_834_data = 32'h0;
  assign RAM_MPORT_834_addr = 10'h342;
  assign RAM_MPORT_834_mask = 1'h1;
  assign RAM_MPORT_834_en = reset;
  assign RAM_MPORT_835_data = 32'h0;
  assign RAM_MPORT_835_addr = 10'h343;
  assign RAM_MPORT_835_mask = 1'h1;
  assign RAM_MPORT_835_en = reset;
  assign RAM_MPORT_836_data = 32'h0;
  assign RAM_MPORT_836_addr = 10'h344;
  assign RAM_MPORT_836_mask = 1'h1;
  assign RAM_MPORT_836_en = reset;
  assign RAM_MPORT_837_data = 32'h0;
  assign RAM_MPORT_837_addr = 10'h345;
  assign RAM_MPORT_837_mask = 1'h1;
  assign RAM_MPORT_837_en = reset;
  assign RAM_MPORT_838_data = 32'h0;
  assign RAM_MPORT_838_addr = 10'h346;
  assign RAM_MPORT_838_mask = 1'h1;
  assign RAM_MPORT_838_en = reset;
  assign RAM_MPORT_839_data = 32'h0;
  assign RAM_MPORT_839_addr = 10'h347;
  assign RAM_MPORT_839_mask = 1'h1;
  assign RAM_MPORT_839_en = reset;
  assign RAM_MPORT_840_data = 32'h0;
  assign RAM_MPORT_840_addr = 10'h348;
  assign RAM_MPORT_840_mask = 1'h1;
  assign RAM_MPORT_840_en = reset;
  assign RAM_MPORT_841_data = 32'h0;
  assign RAM_MPORT_841_addr = 10'h349;
  assign RAM_MPORT_841_mask = 1'h1;
  assign RAM_MPORT_841_en = reset;
  assign RAM_MPORT_842_data = 32'h0;
  assign RAM_MPORT_842_addr = 10'h34a;
  assign RAM_MPORT_842_mask = 1'h1;
  assign RAM_MPORT_842_en = reset;
  assign RAM_MPORT_843_data = 32'h0;
  assign RAM_MPORT_843_addr = 10'h34b;
  assign RAM_MPORT_843_mask = 1'h1;
  assign RAM_MPORT_843_en = reset;
  assign RAM_MPORT_844_data = 32'h0;
  assign RAM_MPORT_844_addr = 10'h34c;
  assign RAM_MPORT_844_mask = 1'h1;
  assign RAM_MPORT_844_en = reset;
  assign RAM_MPORT_845_data = 32'h0;
  assign RAM_MPORT_845_addr = 10'h34d;
  assign RAM_MPORT_845_mask = 1'h1;
  assign RAM_MPORT_845_en = reset;
  assign RAM_MPORT_846_data = 32'h0;
  assign RAM_MPORT_846_addr = 10'h34e;
  assign RAM_MPORT_846_mask = 1'h1;
  assign RAM_MPORT_846_en = reset;
  assign RAM_MPORT_847_data = 32'h0;
  assign RAM_MPORT_847_addr = 10'h34f;
  assign RAM_MPORT_847_mask = 1'h1;
  assign RAM_MPORT_847_en = reset;
  assign RAM_MPORT_848_data = 32'h0;
  assign RAM_MPORT_848_addr = 10'h350;
  assign RAM_MPORT_848_mask = 1'h1;
  assign RAM_MPORT_848_en = reset;
  assign RAM_MPORT_849_data = 32'h0;
  assign RAM_MPORT_849_addr = 10'h351;
  assign RAM_MPORT_849_mask = 1'h1;
  assign RAM_MPORT_849_en = reset;
  assign RAM_MPORT_850_data = 32'h0;
  assign RAM_MPORT_850_addr = 10'h352;
  assign RAM_MPORT_850_mask = 1'h1;
  assign RAM_MPORT_850_en = reset;
  assign RAM_MPORT_851_data = 32'h0;
  assign RAM_MPORT_851_addr = 10'h353;
  assign RAM_MPORT_851_mask = 1'h1;
  assign RAM_MPORT_851_en = reset;
  assign RAM_MPORT_852_data = 32'h0;
  assign RAM_MPORT_852_addr = 10'h354;
  assign RAM_MPORT_852_mask = 1'h1;
  assign RAM_MPORT_852_en = reset;
  assign RAM_MPORT_853_data = 32'h0;
  assign RAM_MPORT_853_addr = 10'h355;
  assign RAM_MPORT_853_mask = 1'h1;
  assign RAM_MPORT_853_en = reset;
  assign RAM_MPORT_854_data = 32'h0;
  assign RAM_MPORT_854_addr = 10'h356;
  assign RAM_MPORT_854_mask = 1'h1;
  assign RAM_MPORT_854_en = reset;
  assign RAM_MPORT_855_data = 32'h0;
  assign RAM_MPORT_855_addr = 10'h357;
  assign RAM_MPORT_855_mask = 1'h1;
  assign RAM_MPORT_855_en = reset;
  assign RAM_MPORT_856_data = 32'h0;
  assign RAM_MPORT_856_addr = 10'h358;
  assign RAM_MPORT_856_mask = 1'h1;
  assign RAM_MPORT_856_en = reset;
  assign RAM_MPORT_857_data = 32'h0;
  assign RAM_MPORT_857_addr = 10'h359;
  assign RAM_MPORT_857_mask = 1'h1;
  assign RAM_MPORT_857_en = reset;
  assign RAM_MPORT_858_data = 32'h0;
  assign RAM_MPORT_858_addr = 10'h35a;
  assign RAM_MPORT_858_mask = 1'h1;
  assign RAM_MPORT_858_en = reset;
  assign RAM_MPORT_859_data = 32'h0;
  assign RAM_MPORT_859_addr = 10'h35b;
  assign RAM_MPORT_859_mask = 1'h1;
  assign RAM_MPORT_859_en = reset;
  assign RAM_MPORT_860_data = 32'h0;
  assign RAM_MPORT_860_addr = 10'h35c;
  assign RAM_MPORT_860_mask = 1'h1;
  assign RAM_MPORT_860_en = reset;
  assign RAM_MPORT_861_data = 32'h0;
  assign RAM_MPORT_861_addr = 10'h35d;
  assign RAM_MPORT_861_mask = 1'h1;
  assign RAM_MPORT_861_en = reset;
  assign RAM_MPORT_862_data = 32'h0;
  assign RAM_MPORT_862_addr = 10'h35e;
  assign RAM_MPORT_862_mask = 1'h1;
  assign RAM_MPORT_862_en = reset;
  assign RAM_MPORT_863_data = 32'h0;
  assign RAM_MPORT_863_addr = 10'h35f;
  assign RAM_MPORT_863_mask = 1'h1;
  assign RAM_MPORT_863_en = reset;
  assign RAM_MPORT_864_data = 32'h0;
  assign RAM_MPORT_864_addr = 10'h360;
  assign RAM_MPORT_864_mask = 1'h1;
  assign RAM_MPORT_864_en = reset;
  assign RAM_MPORT_865_data = 32'h0;
  assign RAM_MPORT_865_addr = 10'h361;
  assign RAM_MPORT_865_mask = 1'h1;
  assign RAM_MPORT_865_en = reset;
  assign RAM_MPORT_866_data = 32'h0;
  assign RAM_MPORT_866_addr = 10'h362;
  assign RAM_MPORT_866_mask = 1'h1;
  assign RAM_MPORT_866_en = reset;
  assign RAM_MPORT_867_data = 32'h0;
  assign RAM_MPORT_867_addr = 10'h363;
  assign RAM_MPORT_867_mask = 1'h1;
  assign RAM_MPORT_867_en = reset;
  assign RAM_MPORT_868_data = 32'h0;
  assign RAM_MPORT_868_addr = 10'h364;
  assign RAM_MPORT_868_mask = 1'h1;
  assign RAM_MPORT_868_en = reset;
  assign RAM_MPORT_869_data = 32'h0;
  assign RAM_MPORT_869_addr = 10'h365;
  assign RAM_MPORT_869_mask = 1'h1;
  assign RAM_MPORT_869_en = reset;
  assign RAM_MPORT_870_data = 32'h0;
  assign RAM_MPORT_870_addr = 10'h366;
  assign RAM_MPORT_870_mask = 1'h1;
  assign RAM_MPORT_870_en = reset;
  assign RAM_MPORT_871_data = 32'h0;
  assign RAM_MPORT_871_addr = 10'h367;
  assign RAM_MPORT_871_mask = 1'h1;
  assign RAM_MPORT_871_en = reset;
  assign RAM_MPORT_872_data = 32'h0;
  assign RAM_MPORT_872_addr = 10'h368;
  assign RAM_MPORT_872_mask = 1'h1;
  assign RAM_MPORT_872_en = reset;
  assign RAM_MPORT_873_data = 32'h0;
  assign RAM_MPORT_873_addr = 10'h369;
  assign RAM_MPORT_873_mask = 1'h1;
  assign RAM_MPORT_873_en = reset;
  assign RAM_MPORT_874_data = 32'h0;
  assign RAM_MPORT_874_addr = 10'h36a;
  assign RAM_MPORT_874_mask = 1'h1;
  assign RAM_MPORT_874_en = reset;
  assign RAM_MPORT_875_data = 32'h0;
  assign RAM_MPORT_875_addr = 10'h36b;
  assign RAM_MPORT_875_mask = 1'h1;
  assign RAM_MPORT_875_en = reset;
  assign RAM_MPORT_876_data = 32'h0;
  assign RAM_MPORT_876_addr = 10'h36c;
  assign RAM_MPORT_876_mask = 1'h1;
  assign RAM_MPORT_876_en = reset;
  assign RAM_MPORT_877_data = 32'h0;
  assign RAM_MPORT_877_addr = 10'h36d;
  assign RAM_MPORT_877_mask = 1'h1;
  assign RAM_MPORT_877_en = reset;
  assign RAM_MPORT_878_data = 32'h0;
  assign RAM_MPORT_878_addr = 10'h36e;
  assign RAM_MPORT_878_mask = 1'h1;
  assign RAM_MPORT_878_en = reset;
  assign RAM_MPORT_879_data = 32'h0;
  assign RAM_MPORT_879_addr = 10'h36f;
  assign RAM_MPORT_879_mask = 1'h1;
  assign RAM_MPORT_879_en = reset;
  assign RAM_MPORT_880_data = 32'h0;
  assign RAM_MPORT_880_addr = 10'h370;
  assign RAM_MPORT_880_mask = 1'h1;
  assign RAM_MPORT_880_en = reset;
  assign RAM_MPORT_881_data = 32'h0;
  assign RAM_MPORT_881_addr = 10'h371;
  assign RAM_MPORT_881_mask = 1'h1;
  assign RAM_MPORT_881_en = reset;
  assign RAM_MPORT_882_data = 32'h0;
  assign RAM_MPORT_882_addr = 10'h372;
  assign RAM_MPORT_882_mask = 1'h1;
  assign RAM_MPORT_882_en = reset;
  assign RAM_MPORT_883_data = 32'h0;
  assign RAM_MPORT_883_addr = 10'h373;
  assign RAM_MPORT_883_mask = 1'h1;
  assign RAM_MPORT_883_en = reset;
  assign RAM_MPORT_884_data = 32'h0;
  assign RAM_MPORT_884_addr = 10'h374;
  assign RAM_MPORT_884_mask = 1'h1;
  assign RAM_MPORT_884_en = reset;
  assign RAM_MPORT_885_data = 32'h0;
  assign RAM_MPORT_885_addr = 10'h375;
  assign RAM_MPORT_885_mask = 1'h1;
  assign RAM_MPORT_885_en = reset;
  assign RAM_MPORT_886_data = 32'h0;
  assign RAM_MPORT_886_addr = 10'h376;
  assign RAM_MPORT_886_mask = 1'h1;
  assign RAM_MPORT_886_en = reset;
  assign RAM_MPORT_887_data = 32'h0;
  assign RAM_MPORT_887_addr = 10'h377;
  assign RAM_MPORT_887_mask = 1'h1;
  assign RAM_MPORT_887_en = reset;
  assign RAM_MPORT_888_data = 32'h0;
  assign RAM_MPORT_888_addr = 10'h378;
  assign RAM_MPORT_888_mask = 1'h1;
  assign RAM_MPORT_888_en = reset;
  assign RAM_MPORT_889_data = 32'h0;
  assign RAM_MPORT_889_addr = 10'h379;
  assign RAM_MPORT_889_mask = 1'h1;
  assign RAM_MPORT_889_en = reset;
  assign RAM_MPORT_890_data = 32'h0;
  assign RAM_MPORT_890_addr = 10'h37a;
  assign RAM_MPORT_890_mask = 1'h1;
  assign RAM_MPORT_890_en = reset;
  assign RAM_MPORT_891_data = 32'h0;
  assign RAM_MPORT_891_addr = 10'h37b;
  assign RAM_MPORT_891_mask = 1'h1;
  assign RAM_MPORT_891_en = reset;
  assign RAM_MPORT_892_data = 32'h0;
  assign RAM_MPORT_892_addr = 10'h37c;
  assign RAM_MPORT_892_mask = 1'h1;
  assign RAM_MPORT_892_en = reset;
  assign RAM_MPORT_893_data = 32'h0;
  assign RAM_MPORT_893_addr = 10'h37d;
  assign RAM_MPORT_893_mask = 1'h1;
  assign RAM_MPORT_893_en = reset;
  assign RAM_MPORT_894_data = 32'h0;
  assign RAM_MPORT_894_addr = 10'h37e;
  assign RAM_MPORT_894_mask = 1'h1;
  assign RAM_MPORT_894_en = reset;
  assign RAM_MPORT_895_data = 32'h0;
  assign RAM_MPORT_895_addr = 10'h37f;
  assign RAM_MPORT_895_mask = 1'h1;
  assign RAM_MPORT_895_en = reset;
  assign RAM_MPORT_896_data = 32'h0;
  assign RAM_MPORT_896_addr = 10'h380;
  assign RAM_MPORT_896_mask = 1'h1;
  assign RAM_MPORT_896_en = reset;
  assign RAM_MPORT_897_data = 32'h0;
  assign RAM_MPORT_897_addr = 10'h381;
  assign RAM_MPORT_897_mask = 1'h1;
  assign RAM_MPORT_897_en = reset;
  assign RAM_MPORT_898_data = 32'h0;
  assign RAM_MPORT_898_addr = 10'h382;
  assign RAM_MPORT_898_mask = 1'h1;
  assign RAM_MPORT_898_en = reset;
  assign RAM_MPORT_899_data = 32'h0;
  assign RAM_MPORT_899_addr = 10'h383;
  assign RAM_MPORT_899_mask = 1'h1;
  assign RAM_MPORT_899_en = reset;
  assign RAM_MPORT_900_data = 32'h0;
  assign RAM_MPORT_900_addr = 10'h384;
  assign RAM_MPORT_900_mask = 1'h1;
  assign RAM_MPORT_900_en = reset;
  assign RAM_MPORT_901_data = 32'h0;
  assign RAM_MPORT_901_addr = 10'h385;
  assign RAM_MPORT_901_mask = 1'h1;
  assign RAM_MPORT_901_en = reset;
  assign RAM_MPORT_902_data = 32'h0;
  assign RAM_MPORT_902_addr = 10'h386;
  assign RAM_MPORT_902_mask = 1'h1;
  assign RAM_MPORT_902_en = reset;
  assign RAM_MPORT_903_data = 32'h0;
  assign RAM_MPORT_903_addr = 10'h387;
  assign RAM_MPORT_903_mask = 1'h1;
  assign RAM_MPORT_903_en = reset;
  assign RAM_MPORT_904_data = 32'h0;
  assign RAM_MPORT_904_addr = 10'h388;
  assign RAM_MPORT_904_mask = 1'h1;
  assign RAM_MPORT_904_en = reset;
  assign RAM_MPORT_905_data = 32'h0;
  assign RAM_MPORT_905_addr = 10'h389;
  assign RAM_MPORT_905_mask = 1'h1;
  assign RAM_MPORT_905_en = reset;
  assign RAM_MPORT_906_data = 32'h0;
  assign RAM_MPORT_906_addr = 10'h38a;
  assign RAM_MPORT_906_mask = 1'h1;
  assign RAM_MPORT_906_en = reset;
  assign RAM_MPORT_907_data = 32'h0;
  assign RAM_MPORT_907_addr = 10'h38b;
  assign RAM_MPORT_907_mask = 1'h1;
  assign RAM_MPORT_907_en = reset;
  assign RAM_MPORT_908_data = 32'h0;
  assign RAM_MPORT_908_addr = 10'h38c;
  assign RAM_MPORT_908_mask = 1'h1;
  assign RAM_MPORT_908_en = reset;
  assign RAM_MPORT_909_data = 32'h0;
  assign RAM_MPORT_909_addr = 10'h38d;
  assign RAM_MPORT_909_mask = 1'h1;
  assign RAM_MPORT_909_en = reset;
  assign RAM_MPORT_910_data = 32'h0;
  assign RAM_MPORT_910_addr = 10'h38e;
  assign RAM_MPORT_910_mask = 1'h1;
  assign RAM_MPORT_910_en = reset;
  assign RAM_MPORT_911_data = 32'h0;
  assign RAM_MPORT_911_addr = 10'h38f;
  assign RAM_MPORT_911_mask = 1'h1;
  assign RAM_MPORT_911_en = reset;
  assign RAM_MPORT_912_data = 32'h0;
  assign RAM_MPORT_912_addr = 10'h390;
  assign RAM_MPORT_912_mask = 1'h1;
  assign RAM_MPORT_912_en = reset;
  assign RAM_MPORT_913_data = 32'h0;
  assign RAM_MPORT_913_addr = 10'h391;
  assign RAM_MPORT_913_mask = 1'h1;
  assign RAM_MPORT_913_en = reset;
  assign RAM_MPORT_914_data = 32'h0;
  assign RAM_MPORT_914_addr = 10'h392;
  assign RAM_MPORT_914_mask = 1'h1;
  assign RAM_MPORT_914_en = reset;
  assign RAM_MPORT_915_data = 32'h0;
  assign RAM_MPORT_915_addr = 10'h393;
  assign RAM_MPORT_915_mask = 1'h1;
  assign RAM_MPORT_915_en = reset;
  assign RAM_MPORT_916_data = 32'h0;
  assign RAM_MPORT_916_addr = 10'h394;
  assign RAM_MPORT_916_mask = 1'h1;
  assign RAM_MPORT_916_en = reset;
  assign RAM_MPORT_917_data = 32'h0;
  assign RAM_MPORT_917_addr = 10'h395;
  assign RAM_MPORT_917_mask = 1'h1;
  assign RAM_MPORT_917_en = reset;
  assign RAM_MPORT_918_data = 32'h0;
  assign RAM_MPORT_918_addr = 10'h396;
  assign RAM_MPORT_918_mask = 1'h1;
  assign RAM_MPORT_918_en = reset;
  assign RAM_MPORT_919_data = 32'h0;
  assign RAM_MPORT_919_addr = 10'h397;
  assign RAM_MPORT_919_mask = 1'h1;
  assign RAM_MPORT_919_en = reset;
  assign RAM_MPORT_920_data = 32'h0;
  assign RAM_MPORT_920_addr = 10'h398;
  assign RAM_MPORT_920_mask = 1'h1;
  assign RAM_MPORT_920_en = reset;
  assign RAM_MPORT_921_data = 32'h0;
  assign RAM_MPORT_921_addr = 10'h399;
  assign RAM_MPORT_921_mask = 1'h1;
  assign RAM_MPORT_921_en = reset;
  assign RAM_MPORT_922_data = 32'h0;
  assign RAM_MPORT_922_addr = 10'h39a;
  assign RAM_MPORT_922_mask = 1'h1;
  assign RAM_MPORT_922_en = reset;
  assign RAM_MPORT_923_data = 32'h0;
  assign RAM_MPORT_923_addr = 10'h39b;
  assign RAM_MPORT_923_mask = 1'h1;
  assign RAM_MPORT_923_en = reset;
  assign RAM_MPORT_924_data = 32'h0;
  assign RAM_MPORT_924_addr = 10'h39c;
  assign RAM_MPORT_924_mask = 1'h1;
  assign RAM_MPORT_924_en = reset;
  assign RAM_MPORT_925_data = 32'h0;
  assign RAM_MPORT_925_addr = 10'h39d;
  assign RAM_MPORT_925_mask = 1'h1;
  assign RAM_MPORT_925_en = reset;
  assign RAM_MPORT_926_data = 32'h0;
  assign RAM_MPORT_926_addr = 10'h39e;
  assign RAM_MPORT_926_mask = 1'h1;
  assign RAM_MPORT_926_en = reset;
  assign RAM_MPORT_927_data = 32'h0;
  assign RAM_MPORT_927_addr = 10'h39f;
  assign RAM_MPORT_927_mask = 1'h1;
  assign RAM_MPORT_927_en = reset;
  assign RAM_MPORT_928_data = 32'h0;
  assign RAM_MPORT_928_addr = 10'h3a0;
  assign RAM_MPORT_928_mask = 1'h1;
  assign RAM_MPORT_928_en = reset;
  assign RAM_MPORT_929_data = 32'h0;
  assign RAM_MPORT_929_addr = 10'h3a1;
  assign RAM_MPORT_929_mask = 1'h1;
  assign RAM_MPORT_929_en = reset;
  assign RAM_MPORT_930_data = 32'h0;
  assign RAM_MPORT_930_addr = 10'h3a2;
  assign RAM_MPORT_930_mask = 1'h1;
  assign RAM_MPORT_930_en = reset;
  assign RAM_MPORT_931_data = 32'h0;
  assign RAM_MPORT_931_addr = 10'h3a3;
  assign RAM_MPORT_931_mask = 1'h1;
  assign RAM_MPORT_931_en = reset;
  assign RAM_MPORT_932_data = 32'h0;
  assign RAM_MPORT_932_addr = 10'h3a4;
  assign RAM_MPORT_932_mask = 1'h1;
  assign RAM_MPORT_932_en = reset;
  assign RAM_MPORT_933_data = 32'h0;
  assign RAM_MPORT_933_addr = 10'h3a5;
  assign RAM_MPORT_933_mask = 1'h1;
  assign RAM_MPORT_933_en = reset;
  assign RAM_MPORT_934_data = 32'h0;
  assign RAM_MPORT_934_addr = 10'h3a6;
  assign RAM_MPORT_934_mask = 1'h1;
  assign RAM_MPORT_934_en = reset;
  assign RAM_MPORT_935_data = 32'h0;
  assign RAM_MPORT_935_addr = 10'h3a7;
  assign RAM_MPORT_935_mask = 1'h1;
  assign RAM_MPORT_935_en = reset;
  assign RAM_MPORT_936_data = 32'h0;
  assign RAM_MPORT_936_addr = 10'h3a8;
  assign RAM_MPORT_936_mask = 1'h1;
  assign RAM_MPORT_936_en = reset;
  assign RAM_MPORT_937_data = 32'h0;
  assign RAM_MPORT_937_addr = 10'h3a9;
  assign RAM_MPORT_937_mask = 1'h1;
  assign RAM_MPORT_937_en = reset;
  assign RAM_MPORT_938_data = 32'h0;
  assign RAM_MPORT_938_addr = 10'h3aa;
  assign RAM_MPORT_938_mask = 1'h1;
  assign RAM_MPORT_938_en = reset;
  assign RAM_MPORT_939_data = 32'h0;
  assign RAM_MPORT_939_addr = 10'h3ab;
  assign RAM_MPORT_939_mask = 1'h1;
  assign RAM_MPORT_939_en = reset;
  assign RAM_MPORT_940_data = 32'h0;
  assign RAM_MPORT_940_addr = 10'h3ac;
  assign RAM_MPORT_940_mask = 1'h1;
  assign RAM_MPORT_940_en = reset;
  assign RAM_MPORT_941_data = 32'h0;
  assign RAM_MPORT_941_addr = 10'h3ad;
  assign RAM_MPORT_941_mask = 1'h1;
  assign RAM_MPORT_941_en = reset;
  assign RAM_MPORT_942_data = 32'h0;
  assign RAM_MPORT_942_addr = 10'h3ae;
  assign RAM_MPORT_942_mask = 1'h1;
  assign RAM_MPORT_942_en = reset;
  assign RAM_MPORT_943_data = 32'h0;
  assign RAM_MPORT_943_addr = 10'h3af;
  assign RAM_MPORT_943_mask = 1'h1;
  assign RAM_MPORT_943_en = reset;
  assign RAM_MPORT_944_data = 32'h0;
  assign RAM_MPORT_944_addr = 10'h3b0;
  assign RAM_MPORT_944_mask = 1'h1;
  assign RAM_MPORT_944_en = reset;
  assign RAM_MPORT_945_data = 32'h0;
  assign RAM_MPORT_945_addr = 10'h3b1;
  assign RAM_MPORT_945_mask = 1'h1;
  assign RAM_MPORT_945_en = reset;
  assign RAM_MPORT_946_data = 32'h0;
  assign RAM_MPORT_946_addr = 10'h3b2;
  assign RAM_MPORT_946_mask = 1'h1;
  assign RAM_MPORT_946_en = reset;
  assign RAM_MPORT_947_data = 32'h0;
  assign RAM_MPORT_947_addr = 10'h3b3;
  assign RAM_MPORT_947_mask = 1'h1;
  assign RAM_MPORT_947_en = reset;
  assign RAM_MPORT_948_data = 32'h0;
  assign RAM_MPORT_948_addr = 10'h3b4;
  assign RAM_MPORT_948_mask = 1'h1;
  assign RAM_MPORT_948_en = reset;
  assign RAM_MPORT_949_data = 32'h0;
  assign RAM_MPORT_949_addr = 10'h3b5;
  assign RAM_MPORT_949_mask = 1'h1;
  assign RAM_MPORT_949_en = reset;
  assign RAM_MPORT_950_data = 32'h0;
  assign RAM_MPORT_950_addr = 10'h3b6;
  assign RAM_MPORT_950_mask = 1'h1;
  assign RAM_MPORT_950_en = reset;
  assign RAM_MPORT_951_data = 32'h0;
  assign RAM_MPORT_951_addr = 10'h3b7;
  assign RAM_MPORT_951_mask = 1'h1;
  assign RAM_MPORT_951_en = reset;
  assign RAM_MPORT_952_data = 32'h0;
  assign RAM_MPORT_952_addr = 10'h3b8;
  assign RAM_MPORT_952_mask = 1'h1;
  assign RAM_MPORT_952_en = reset;
  assign RAM_MPORT_953_data = 32'h0;
  assign RAM_MPORT_953_addr = 10'h3b9;
  assign RAM_MPORT_953_mask = 1'h1;
  assign RAM_MPORT_953_en = reset;
  assign RAM_MPORT_954_data = 32'h0;
  assign RAM_MPORT_954_addr = 10'h3ba;
  assign RAM_MPORT_954_mask = 1'h1;
  assign RAM_MPORT_954_en = reset;
  assign RAM_MPORT_955_data = 32'h0;
  assign RAM_MPORT_955_addr = 10'h3bb;
  assign RAM_MPORT_955_mask = 1'h1;
  assign RAM_MPORT_955_en = reset;
  assign RAM_MPORT_956_data = 32'h0;
  assign RAM_MPORT_956_addr = 10'h3bc;
  assign RAM_MPORT_956_mask = 1'h1;
  assign RAM_MPORT_956_en = reset;
  assign RAM_MPORT_957_data = 32'h0;
  assign RAM_MPORT_957_addr = 10'h3bd;
  assign RAM_MPORT_957_mask = 1'h1;
  assign RAM_MPORT_957_en = reset;
  assign RAM_MPORT_958_data = 32'h0;
  assign RAM_MPORT_958_addr = 10'h3be;
  assign RAM_MPORT_958_mask = 1'h1;
  assign RAM_MPORT_958_en = reset;
  assign RAM_MPORT_959_data = 32'h0;
  assign RAM_MPORT_959_addr = 10'h3bf;
  assign RAM_MPORT_959_mask = 1'h1;
  assign RAM_MPORT_959_en = reset;
  assign RAM_MPORT_960_data = 32'h0;
  assign RAM_MPORT_960_addr = 10'h3c0;
  assign RAM_MPORT_960_mask = 1'h1;
  assign RAM_MPORT_960_en = reset;
  assign RAM_MPORT_961_data = 32'h0;
  assign RAM_MPORT_961_addr = 10'h3c1;
  assign RAM_MPORT_961_mask = 1'h1;
  assign RAM_MPORT_961_en = reset;
  assign RAM_MPORT_962_data = 32'h0;
  assign RAM_MPORT_962_addr = 10'h3c2;
  assign RAM_MPORT_962_mask = 1'h1;
  assign RAM_MPORT_962_en = reset;
  assign RAM_MPORT_963_data = 32'h0;
  assign RAM_MPORT_963_addr = 10'h3c3;
  assign RAM_MPORT_963_mask = 1'h1;
  assign RAM_MPORT_963_en = reset;
  assign RAM_MPORT_964_data = 32'h0;
  assign RAM_MPORT_964_addr = 10'h3c4;
  assign RAM_MPORT_964_mask = 1'h1;
  assign RAM_MPORT_964_en = reset;
  assign RAM_MPORT_965_data = 32'h0;
  assign RAM_MPORT_965_addr = 10'h3c5;
  assign RAM_MPORT_965_mask = 1'h1;
  assign RAM_MPORT_965_en = reset;
  assign RAM_MPORT_966_data = 32'h0;
  assign RAM_MPORT_966_addr = 10'h3c6;
  assign RAM_MPORT_966_mask = 1'h1;
  assign RAM_MPORT_966_en = reset;
  assign RAM_MPORT_967_data = 32'h0;
  assign RAM_MPORT_967_addr = 10'h3c7;
  assign RAM_MPORT_967_mask = 1'h1;
  assign RAM_MPORT_967_en = reset;
  assign RAM_MPORT_968_data = 32'h0;
  assign RAM_MPORT_968_addr = 10'h3c8;
  assign RAM_MPORT_968_mask = 1'h1;
  assign RAM_MPORT_968_en = reset;
  assign RAM_MPORT_969_data = 32'h0;
  assign RAM_MPORT_969_addr = 10'h3c9;
  assign RAM_MPORT_969_mask = 1'h1;
  assign RAM_MPORT_969_en = reset;
  assign RAM_MPORT_970_data = 32'h0;
  assign RAM_MPORT_970_addr = 10'h3ca;
  assign RAM_MPORT_970_mask = 1'h1;
  assign RAM_MPORT_970_en = reset;
  assign RAM_MPORT_971_data = 32'h0;
  assign RAM_MPORT_971_addr = 10'h3cb;
  assign RAM_MPORT_971_mask = 1'h1;
  assign RAM_MPORT_971_en = reset;
  assign RAM_MPORT_972_data = 32'h0;
  assign RAM_MPORT_972_addr = 10'h3cc;
  assign RAM_MPORT_972_mask = 1'h1;
  assign RAM_MPORT_972_en = reset;
  assign RAM_MPORT_973_data = 32'h0;
  assign RAM_MPORT_973_addr = 10'h3cd;
  assign RAM_MPORT_973_mask = 1'h1;
  assign RAM_MPORT_973_en = reset;
  assign RAM_MPORT_974_data = 32'h0;
  assign RAM_MPORT_974_addr = 10'h3ce;
  assign RAM_MPORT_974_mask = 1'h1;
  assign RAM_MPORT_974_en = reset;
  assign RAM_MPORT_975_data = 32'h0;
  assign RAM_MPORT_975_addr = 10'h3cf;
  assign RAM_MPORT_975_mask = 1'h1;
  assign RAM_MPORT_975_en = reset;
  assign RAM_MPORT_976_data = 32'h0;
  assign RAM_MPORT_976_addr = 10'h3d0;
  assign RAM_MPORT_976_mask = 1'h1;
  assign RAM_MPORT_976_en = reset;
  assign RAM_MPORT_977_data = 32'h0;
  assign RAM_MPORT_977_addr = 10'h3d1;
  assign RAM_MPORT_977_mask = 1'h1;
  assign RAM_MPORT_977_en = reset;
  assign RAM_MPORT_978_data = 32'h0;
  assign RAM_MPORT_978_addr = 10'h3d2;
  assign RAM_MPORT_978_mask = 1'h1;
  assign RAM_MPORT_978_en = reset;
  assign RAM_MPORT_979_data = 32'h0;
  assign RAM_MPORT_979_addr = 10'h3d3;
  assign RAM_MPORT_979_mask = 1'h1;
  assign RAM_MPORT_979_en = reset;
  assign RAM_MPORT_980_data = 32'h0;
  assign RAM_MPORT_980_addr = 10'h3d4;
  assign RAM_MPORT_980_mask = 1'h1;
  assign RAM_MPORT_980_en = reset;
  assign RAM_MPORT_981_data = 32'h0;
  assign RAM_MPORT_981_addr = 10'h3d5;
  assign RAM_MPORT_981_mask = 1'h1;
  assign RAM_MPORT_981_en = reset;
  assign RAM_MPORT_982_data = 32'h0;
  assign RAM_MPORT_982_addr = 10'h3d6;
  assign RAM_MPORT_982_mask = 1'h1;
  assign RAM_MPORT_982_en = reset;
  assign RAM_MPORT_983_data = 32'h0;
  assign RAM_MPORT_983_addr = 10'h3d7;
  assign RAM_MPORT_983_mask = 1'h1;
  assign RAM_MPORT_983_en = reset;
  assign RAM_MPORT_984_data = 32'h0;
  assign RAM_MPORT_984_addr = 10'h3d8;
  assign RAM_MPORT_984_mask = 1'h1;
  assign RAM_MPORT_984_en = reset;
  assign RAM_MPORT_985_data = 32'h0;
  assign RAM_MPORT_985_addr = 10'h3d9;
  assign RAM_MPORT_985_mask = 1'h1;
  assign RAM_MPORT_985_en = reset;
  assign RAM_MPORT_986_data = 32'h0;
  assign RAM_MPORT_986_addr = 10'h3da;
  assign RAM_MPORT_986_mask = 1'h1;
  assign RAM_MPORT_986_en = reset;
  assign RAM_MPORT_987_data = 32'h0;
  assign RAM_MPORT_987_addr = 10'h3db;
  assign RAM_MPORT_987_mask = 1'h1;
  assign RAM_MPORT_987_en = reset;
  assign RAM_MPORT_988_data = 32'h0;
  assign RAM_MPORT_988_addr = 10'h3dc;
  assign RAM_MPORT_988_mask = 1'h1;
  assign RAM_MPORT_988_en = reset;
  assign RAM_MPORT_989_data = 32'h0;
  assign RAM_MPORT_989_addr = 10'h3dd;
  assign RAM_MPORT_989_mask = 1'h1;
  assign RAM_MPORT_989_en = reset;
  assign RAM_MPORT_990_data = 32'h0;
  assign RAM_MPORT_990_addr = 10'h3de;
  assign RAM_MPORT_990_mask = 1'h1;
  assign RAM_MPORT_990_en = reset;
  assign RAM_MPORT_991_data = 32'h0;
  assign RAM_MPORT_991_addr = 10'h3df;
  assign RAM_MPORT_991_mask = 1'h1;
  assign RAM_MPORT_991_en = reset;
  assign RAM_MPORT_992_data = 32'h0;
  assign RAM_MPORT_992_addr = 10'h3e0;
  assign RAM_MPORT_992_mask = 1'h1;
  assign RAM_MPORT_992_en = reset;
  assign RAM_MPORT_993_data = 32'h0;
  assign RAM_MPORT_993_addr = 10'h3e1;
  assign RAM_MPORT_993_mask = 1'h1;
  assign RAM_MPORT_993_en = reset;
  assign RAM_MPORT_994_data = 32'h0;
  assign RAM_MPORT_994_addr = 10'h3e2;
  assign RAM_MPORT_994_mask = 1'h1;
  assign RAM_MPORT_994_en = reset;
  assign RAM_MPORT_995_data = 32'h0;
  assign RAM_MPORT_995_addr = 10'h3e3;
  assign RAM_MPORT_995_mask = 1'h1;
  assign RAM_MPORT_995_en = reset;
  assign RAM_MPORT_996_data = 32'h0;
  assign RAM_MPORT_996_addr = 10'h3e4;
  assign RAM_MPORT_996_mask = 1'h1;
  assign RAM_MPORT_996_en = reset;
  assign RAM_MPORT_997_data = 32'h0;
  assign RAM_MPORT_997_addr = 10'h3e5;
  assign RAM_MPORT_997_mask = 1'h1;
  assign RAM_MPORT_997_en = reset;
  assign RAM_MPORT_998_data = 32'h0;
  assign RAM_MPORT_998_addr = 10'h3e6;
  assign RAM_MPORT_998_mask = 1'h1;
  assign RAM_MPORT_998_en = reset;
  assign RAM_MPORT_999_data = 32'h0;
  assign RAM_MPORT_999_addr = 10'h3e7;
  assign RAM_MPORT_999_mask = 1'h1;
  assign RAM_MPORT_999_en = reset;
  assign RAM_MPORT_1000_data = 32'h0;
  assign RAM_MPORT_1000_addr = 10'h3e8;
  assign RAM_MPORT_1000_mask = 1'h1;
  assign RAM_MPORT_1000_en = reset;
  assign RAM_MPORT_1001_data = 32'h0;
  assign RAM_MPORT_1001_addr = 10'h3e9;
  assign RAM_MPORT_1001_mask = 1'h1;
  assign RAM_MPORT_1001_en = reset;
  assign RAM_MPORT_1002_data = 32'h0;
  assign RAM_MPORT_1002_addr = 10'h3ea;
  assign RAM_MPORT_1002_mask = 1'h1;
  assign RAM_MPORT_1002_en = reset;
  assign RAM_MPORT_1003_data = 32'h0;
  assign RAM_MPORT_1003_addr = 10'h3eb;
  assign RAM_MPORT_1003_mask = 1'h1;
  assign RAM_MPORT_1003_en = reset;
  assign RAM_MPORT_1004_data = 32'h0;
  assign RAM_MPORT_1004_addr = 10'h3ec;
  assign RAM_MPORT_1004_mask = 1'h1;
  assign RAM_MPORT_1004_en = reset;
  assign RAM_MPORT_1005_data = 32'h0;
  assign RAM_MPORT_1005_addr = 10'h3ed;
  assign RAM_MPORT_1005_mask = 1'h1;
  assign RAM_MPORT_1005_en = reset;
  assign RAM_MPORT_1006_data = 32'h0;
  assign RAM_MPORT_1006_addr = 10'h3ee;
  assign RAM_MPORT_1006_mask = 1'h1;
  assign RAM_MPORT_1006_en = reset;
  assign RAM_MPORT_1007_data = 32'h0;
  assign RAM_MPORT_1007_addr = 10'h3ef;
  assign RAM_MPORT_1007_mask = 1'h1;
  assign RAM_MPORT_1007_en = reset;
  assign RAM_MPORT_1008_data = 32'h0;
  assign RAM_MPORT_1008_addr = 10'h3f0;
  assign RAM_MPORT_1008_mask = 1'h1;
  assign RAM_MPORT_1008_en = reset;
  assign RAM_MPORT_1009_data = 32'h0;
  assign RAM_MPORT_1009_addr = 10'h3f1;
  assign RAM_MPORT_1009_mask = 1'h1;
  assign RAM_MPORT_1009_en = reset;
  assign RAM_MPORT_1010_data = 32'h0;
  assign RAM_MPORT_1010_addr = 10'h3f2;
  assign RAM_MPORT_1010_mask = 1'h1;
  assign RAM_MPORT_1010_en = reset;
  assign RAM_MPORT_1011_data = 32'h0;
  assign RAM_MPORT_1011_addr = 10'h3f3;
  assign RAM_MPORT_1011_mask = 1'h1;
  assign RAM_MPORT_1011_en = reset;
  assign RAM_MPORT_1012_data = 32'h0;
  assign RAM_MPORT_1012_addr = 10'h3f4;
  assign RAM_MPORT_1012_mask = 1'h1;
  assign RAM_MPORT_1012_en = reset;
  assign RAM_MPORT_1013_data = 32'h0;
  assign RAM_MPORT_1013_addr = 10'h3f5;
  assign RAM_MPORT_1013_mask = 1'h1;
  assign RAM_MPORT_1013_en = reset;
  assign RAM_MPORT_1014_data = 32'h0;
  assign RAM_MPORT_1014_addr = 10'h3f6;
  assign RAM_MPORT_1014_mask = 1'h1;
  assign RAM_MPORT_1014_en = reset;
  assign RAM_MPORT_1015_data = 32'h0;
  assign RAM_MPORT_1015_addr = 10'h3f7;
  assign RAM_MPORT_1015_mask = 1'h1;
  assign RAM_MPORT_1015_en = reset;
  assign RAM_MPORT_1016_data = 32'h0;
  assign RAM_MPORT_1016_addr = 10'h3f8;
  assign RAM_MPORT_1016_mask = 1'h1;
  assign RAM_MPORT_1016_en = reset;
  assign RAM_MPORT_1017_data = 32'h0;
  assign RAM_MPORT_1017_addr = 10'h3f9;
  assign RAM_MPORT_1017_mask = 1'h1;
  assign RAM_MPORT_1017_en = reset;
  assign RAM_MPORT_1018_data = 32'h0;
  assign RAM_MPORT_1018_addr = 10'h3fa;
  assign RAM_MPORT_1018_mask = 1'h1;
  assign RAM_MPORT_1018_en = reset;
  assign RAM_MPORT_1019_data = 32'h0;
  assign RAM_MPORT_1019_addr = 10'h3fb;
  assign RAM_MPORT_1019_mask = 1'h1;
  assign RAM_MPORT_1019_en = reset;
  assign RAM_MPORT_1020_data = 32'h0;
  assign RAM_MPORT_1020_addr = 10'h3fc;
  assign RAM_MPORT_1020_mask = 1'h1;
  assign RAM_MPORT_1020_en = reset;
  assign RAM_MPORT_1021_data = 32'h0;
  assign RAM_MPORT_1021_addr = 10'h3fd;
  assign RAM_MPORT_1021_mask = 1'h1;
  assign RAM_MPORT_1021_en = reset;
  assign RAM_MPORT_1022_data = 32'h0;
  assign RAM_MPORT_1022_addr = 10'h3fe;
  assign RAM_MPORT_1022_mask = 1'h1;
  assign RAM_MPORT_1022_en = reset;
  assign RAM_MPORT_1023_data = 32'h0;
  assign RAM_MPORT_1023_addr = 10'h3ff;
  assign RAM_MPORT_1023_mask = 1'h1;
  assign RAM_MPORT_1023_en = reset;
  assign RAM_MPORT_1024_data = io_WD;
  assign RAM_MPORT_1024_addr = io_Addr[11:2];
  assign RAM_MPORT_1024_mask = 1'h1;
  assign RAM_MPORT_1024_en = reset ? 1'h0 : io_WE;
  assign io_RD = RAM_io_RD_MPORT_data; // @[DM.scala 23:11]
  always @(posedge clock) begin
    if (RAM_MPORT_en & RAM_MPORT_mask) begin
      RAM[RAM_MPORT_addr] <= RAM_MPORT_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1_en & RAM_MPORT_1_mask) begin
      RAM[RAM_MPORT_1_addr] <= RAM_MPORT_1_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_2_en & RAM_MPORT_2_mask) begin
      RAM[RAM_MPORT_2_addr] <= RAM_MPORT_2_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_3_en & RAM_MPORT_3_mask) begin
      RAM[RAM_MPORT_3_addr] <= RAM_MPORT_3_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_4_en & RAM_MPORT_4_mask) begin
      RAM[RAM_MPORT_4_addr] <= RAM_MPORT_4_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_5_en & RAM_MPORT_5_mask) begin
      RAM[RAM_MPORT_5_addr] <= RAM_MPORT_5_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_6_en & RAM_MPORT_6_mask) begin
      RAM[RAM_MPORT_6_addr] <= RAM_MPORT_6_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_7_en & RAM_MPORT_7_mask) begin
      RAM[RAM_MPORT_7_addr] <= RAM_MPORT_7_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_8_en & RAM_MPORT_8_mask) begin
      RAM[RAM_MPORT_8_addr] <= RAM_MPORT_8_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_9_en & RAM_MPORT_9_mask) begin
      RAM[RAM_MPORT_9_addr] <= RAM_MPORT_9_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_10_en & RAM_MPORT_10_mask) begin
      RAM[RAM_MPORT_10_addr] <= RAM_MPORT_10_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_11_en & RAM_MPORT_11_mask) begin
      RAM[RAM_MPORT_11_addr] <= RAM_MPORT_11_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_12_en & RAM_MPORT_12_mask) begin
      RAM[RAM_MPORT_12_addr] <= RAM_MPORT_12_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_13_en & RAM_MPORT_13_mask) begin
      RAM[RAM_MPORT_13_addr] <= RAM_MPORT_13_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_14_en & RAM_MPORT_14_mask) begin
      RAM[RAM_MPORT_14_addr] <= RAM_MPORT_14_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_15_en & RAM_MPORT_15_mask) begin
      RAM[RAM_MPORT_15_addr] <= RAM_MPORT_15_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_16_en & RAM_MPORT_16_mask) begin
      RAM[RAM_MPORT_16_addr] <= RAM_MPORT_16_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_17_en & RAM_MPORT_17_mask) begin
      RAM[RAM_MPORT_17_addr] <= RAM_MPORT_17_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_18_en & RAM_MPORT_18_mask) begin
      RAM[RAM_MPORT_18_addr] <= RAM_MPORT_18_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_19_en & RAM_MPORT_19_mask) begin
      RAM[RAM_MPORT_19_addr] <= RAM_MPORT_19_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_20_en & RAM_MPORT_20_mask) begin
      RAM[RAM_MPORT_20_addr] <= RAM_MPORT_20_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_21_en & RAM_MPORT_21_mask) begin
      RAM[RAM_MPORT_21_addr] <= RAM_MPORT_21_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_22_en & RAM_MPORT_22_mask) begin
      RAM[RAM_MPORT_22_addr] <= RAM_MPORT_22_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_23_en & RAM_MPORT_23_mask) begin
      RAM[RAM_MPORT_23_addr] <= RAM_MPORT_23_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_24_en & RAM_MPORT_24_mask) begin
      RAM[RAM_MPORT_24_addr] <= RAM_MPORT_24_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_25_en & RAM_MPORT_25_mask) begin
      RAM[RAM_MPORT_25_addr] <= RAM_MPORT_25_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_26_en & RAM_MPORT_26_mask) begin
      RAM[RAM_MPORT_26_addr] <= RAM_MPORT_26_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_27_en & RAM_MPORT_27_mask) begin
      RAM[RAM_MPORT_27_addr] <= RAM_MPORT_27_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_28_en & RAM_MPORT_28_mask) begin
      RAM[RAM_MPORT_28_addr] <= RAM_MPORT_28_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_29_en & RAM_MPORT_29_mask) begin
      RAM[RAM_MPORT_29_addr] <= RAM_MPORT_29_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_30_en & RAM_MPORT_30_mask) begin
      RAM[RAM_MPORT_30_addr] <= RAM_MPORT_30_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_31_en & RAM_MPORT_31_mask) begin
      RAM[RAM_MPORT_31_addr] <= RAM_MPORT_31_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_32_en & RAM_MPORT_32_mask) begin
      RAM[RAM_MPORT_32_addr] <= RAM_MPORT_32_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_33_en & RAM_MPORT_33_mask) begin
      RAM[RAM_MPORT_33_addr] <= RAM_MPORT_33_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_34_en & RAM_MPORT_34_mask) begin
      RAM[RAM_MPORT_34_addr] <= RAM_MPORT_34_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_35_en & RAM_MPORT_35_mask) begin
      RAM[RAM_MPORT_35_addr] <= RAM_MPORT_35_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_36_en & RAM_MPORT_36_mask) begin
      RAM[RAM_MPORT_36_addr] <= RAM_MPORT_36_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_37_en & RAM_MPORT_37_mask) begin
      RAM[RAM_MPORT_37_addr] <= RAM_MPORT_37_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_38_en & RAM_MPORT_38_mask) begin
      RAM[RAM_MPORT_38_addr] <= RAM_MPORT_38_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_39_en & RAM_MPORT_39_mask) begin
      RAM[RAM_MPORT_39_addr] <= RAM_MPORT_39_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_40_en & RAM_MPORT_40_mask) begin
      RAM[RAM_MPORT_40_addr] <= RAM_MPORT_40_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_41_en & RAM_MPORT_41_mask) begin
      RAM[RAM_MPORT_41_addr] <= RAM_MPORT_41_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_42_en & RAM_MPORT_42_mask) begin
      RAM[RAM_MPORT_42_addr] <= RAM_MPORT_42_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_43_en & RAM_MPORT_43_mask) begin
      RAM[RAM_MPORT_43_addr] <= RAM_MPORT_43_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_44_en & RAM_MPORT_44_mask) begin
      RAM[RAM_MPORT_44_addr] <= RAM_MPORT_44_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_45_en & RAM_MPORT_45_mask) begin
      RAM[RAM_MPORT_45_addr] <= RAM_MPORT_45_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_46_en & RAM_MPORT_46_mask) begin
      RAM[RAM_MPORT_46_addr] <= RAM_MPORT_46_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_47_en & RAM_MPORT_47_mask) begin
      RAM[RAM_MPORT_47_addr] <= RAM_MPORT_47_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_48_en & RAM_MPORT_48_mask) begin
      RAM[RAM_MPORT_48_addr] <= RAM_MPORT_48_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_49_en & RAM_MPORT_49_mask) begin
      RAM[RAM_MPORT_49_addr] <= RAM_MPORT_49_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_50_en & RAM_MPORT_50_mask) begin
      RAM[RAM_MPORT_50_addr] <= RAM_MPORT_50_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_51_en & RAM_MPORT_51_mask) begin
      RAM[RAM_MPORT_51_addr] <= RAM_MPORT_51_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_52_en & RAM_MPORT_52_mask) begin
      RAM[RAM_MPORT_52_addr] <= RAM_MPORT_52_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_53_en & RAM_MPORT_53_mask) begin
      RAM[RAM_MPORT_53_addr] <= RAM_MPORT_53_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_54_en & RAM_MPORT_54_mask) begin
      RAM[RAM_MPORT_54_addr] <= RAM_MPORT_54_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_55_en & RAM_MPORT_55_mask) begin
      RAM[RAM_MPORT_55_addr] <= RAM_MPORT_55_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_56_en & RAM_MPORT_56_mask) begin
      RAM[RAM_MPORT_56_addr] <= RAM_MPORT_56_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_57_en & RAM_MPORT_57_mask) begin
      RAM[RAM_MPORT_57_addr] <= RAM_MPORT_57_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_58_en & RAM_MPORT_58_mask) begin
      RAM[RAM_MPORT_58_addr] <= RAM_MPORT_58_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_59_en & RAM_MPORT_59_mask) begin
      RAM[RAM_MPORT_59_addr] <= RAM_MPORT_59_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_60_en & RAM_MPORT_60_mask) begin
      RAM[RAM_MPORT_60_addr] <= RAM_MPORT_60_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_61_en & RAM_MPORT_61_mask) begin
      RAM[RAM_MPORT_61_addr] <= RAM_MPORT_61_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_62_en & RAM_MPORT_62_mask) begin
      RAM[RAM_MPORT_62_addr] <= RAM_MPORT_62_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_63_en & RAM_MPORT_63_mask) begin
      RAM[RAM_MPORT_63_addr] <= RAM_MPORT_63_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_64_en & RAM_MPORT_64_mask) begin
      RAM[RAM_MPORT_64_addr] <= RAM_MPORT_64_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_65_en & RAM_MPORT_65_mask) begin
      RAM[RAM_MPORT_65_addr] <= RAM_MPORT_65_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_66_en & RAM_MPORT_66_mask) begin
      RAM[RAM_MPORT_66_addr] <= RAM_MPORT_66_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_67_en & RAM_MPORT_67_mask) begin
      RAM[RAM_MPORT_67_addr] <= RAM_MPORT_67_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_68_en & RAM_MPORT_68_mask) begin
      RAM[RAM_MPORT_68_addr] <= RAM_MPORT_68_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_69_en & RAM_MPORT_69_mask) begin
      RAM[RAM_MPORT_69_addr] <= RAM_MPORT_69_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_70_en & RAM_MPORT_70_mask) begin
      RAM[RAM_MPORT_70_addr] <= RAM_MPORT_70_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_71_en & RAM_MPORT_71_mask) begin
      RAM[RAM_MPORT_71_addr] <= RAM_MPORT_71_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_72_en & RAM_MPORT_72_mask) begin
      RAM[RAM_MPORT_72_addr] <= RAM_MPORT_72_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_73_en & RAM_MPORT_73_mask) begin
      RAM[RAM_MPORT_73_addr] <= RAM_MPORT_73_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_74_en & RAM_MPORT_74_mask) begin
      RAM[RAM_MPORT_74_addr] <= RAM_MPORT_74_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_75_en & RAM_MPORT_75_mask) begin
      RAM[RAM_MPORT_75_addr] <= RAM_MPORT_75_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_76_en & RAM_MPORT_76_mask) begin
      RAM[RAM_MPORT_76_addr] <= RAM_MPORT_76_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_77_en & RAM_MPORT_77_mask) begin
      RAM[RAM_MPORT_77_addr] <= RAM_MPORT_77_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_78_en & RAM_MPORT_78_mask) begin
      RAM[RAM_MPORT_78_addr] <= RAM_MPORT_78_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_79_en & RAM_MPORT_79_mask) begin
      RAM[RAM_MPORT_79_addr] <= RAM_MPORT_79_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_80_en & RAM_MPORT_80_mask) begin
      RAM[RAM_MPORT_80_addr] <= RAM_MPORT_80_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_81_en & RAM_MPORT_81_mask) begin
      RAM[RAM_MPORT_81_addr] <= RAM_MPORT_81_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_82_en & RAM_MPORT_82_mask) begin
      RAM[RAM_MPORT_82_addr] <= RAM_MPORT_82_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_83_en & RAM_MPORT_83_mask) begin
      RAM[RAM_MPORT_83_addr] <= RAM_MPORT_83_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_84_en & RAM_MPORT_84_mask) begin
      RAM[RAM_MPORT_84_addr] <= RAM_MPORT_84_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_85_en & RAM_MPORT_85_mask) begin
      RAM[RAM_MPORT_85_addr] <= RAM_MPORT_85_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_86_en & RAM_MPORT_86_mask) begin
      RAM[RAM_MPORT_86_addr] <= RAM_MPORT_86_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_87_en & RAM_MPORT_87_mask) begin
      RAM[RAM_MPORT_87_addr] <= RAM_MPORT_87_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_88_en & RAM_MPORT_88_mask) begin
      RAM[RAM_MPORT_88_addr] <= RAM_MPORT_88_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_89_en & RAM_MPORT_89_mask) begin
      RAM[RAM_MPORT_89_addr] <= RAM_MPORT_89_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_90_en & RAM_MPORT_90_mask) begin
      RAM[RAM_MPORT_90_addr] <= RAM_MPORT_90_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_91_en & RAM_MPORT_91_mask) begin
      RAM[RAM_MPORT_91_addr] <= RAM_MPORT_91_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_92_en & RAM_MPORT_92_mask) begin
      RAM[RAM_MPORT_92_addr] <= RAM_MPORT_92_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_93_en & RAM_MPORT_93_mask) begin
      RAM[RAM_MPORT_93_addr] <= RAM_MPORT_93_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_94_en & RAM_MPORT_94_mask) begin
      RAM[RAM_MPORT_94_addr] <= RAM_MPORT_94_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_95_en & RAM_MPORT_95_mask) begin
      RAM[RAM_MPORT_95_addr] <= RAM_MPORT_95_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_96_en & RAM_MPORT_96_mask) begin
      RAM[RAM_MPORT_96_addr] <= RAM_MPORT_96_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_97_en & RAM_MPORT_97_mask) begin
      RAM[RAM_MPORT_97_addr] <= RAM_MPORT_97_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_98_en & RAM_MPORT_98_mask) begin
      RAM[RAM_MPORT_98_addr] <= RAM_MPORT_98_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_99_en & RAM_MPORT_99_mask) begin
      RAM[RAM_MPORT_99_addr] <= RAM_MPORT_99_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_100_en & RAM_MPORT_100_mask) begin
      RAM[RAM_MPORT_100_addr] <= RAM_MPORT_100_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_101_en & RAM_MPORT_101_mask) begin
      RAM[RAM_MPORT_101_addr] <= RAM_MPORT_101_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_102_en & RAM_MPORT_102_mask) begin
      RAM[RAM_MPORT_102_addr] <= RAM_MPORT_102_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_103_en & RAM_MPORT_103_mask) begin
      RAM[RAM_MPORT_103_addr] <= RAM_MPORT_103_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_104_en & RAM_MPORT_104_mask) begin
      RAM[RAM_MPORT_104_addr] <= RAM_MPORT_104_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_105_en & RAM_MPORT_105_mask) begin
      RAM[RAM_MPORT_105_addr] <= RAM_MPORT_105_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_106_en & RAM_MPORT_106_mask) begin
      RAM[RAM_MPORT_106_addr] <= RAM_MPORT_106_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_107_en & RAM_MPORT_107_mask) begin
      RAM[RAM_MPORT_107_addr] <= RAM_MPORT_107_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_108_en & RAM_MPORT_108_mask) begin
      RAM[RAM_MPORT_108_addr] <= RAM_MPORT_108_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_109_en & RAM_MPORT_109_mask) begin
      RAM[RAM_MPORT_109_addr] <= RAM_MPORT_109_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_110_en & RAM_MPORT_110_mask) begin
      RAM[RAM_MPORT_110_addr] <= RAM_MPORT_110_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_111_en & RAM_MPORT_111_mask) begin
      RAM[RAM_MPORT_111_addr] <= RAM_MPORT_111_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_112_en & RAM_MPORT_112_mask) begin
      RAM[RAM_MPORT_112_addr] <= RAM_MPORT_112_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_113_en & RAM_MPORT_113_mask) begin
      RAM[RAM_MPORT_113_addr] <= RAM_MPORT_113_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_114_en & RAM_MPORT_114_mask) begin
      RAM[RAM_MPORT_114_addr] <= RAM_MPORT_114_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_115_en & RAM_MPORT_115_mask) begin
      RAM[RAM_MPORT_115_addr] <= RAM_MPORT_115_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_116_en & RAM_MPORT_116_mask) begin
      RAM[RAM_MPORT_116_addr] <= RAM_MPORT_116_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_117_en & RAM_MPORT_117_mask) begin
      RAM[RAM_MPORT_117_addr] <= RAM_MPORT_117_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_118_en & RAM_MPORT_118_mask) begin
      RAM[RAM_MPORT_118_addr] <= RAM_MPORT_118_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_119_en & RAM_MPORT_119_mask) begin
      RAM[RAM_MPORT_119_addr] <= RAM_MPORT_119_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_120_en & RAM_MPORT_120_mask) begin
      RAM[RAM_MPORT_120_addr] <= RAM_MPORT_120_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_121_en & RAM_MPORT_121_mask) begin
      RAM[RAM_MPORT_121_addr] <= RAM_MPORT_121_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_122_en & RAM_MPORT_122_mask) begin
      RAM[RAM_MPORT_122_addr] <= RAM_MPORT_122_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_123_en & RAM_MPORT_123_mask) begin
      RAM[RAM_MPORT_123_addr] <= RAM_MPORT_123_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_124_en & RAM_MPORT_124_mask) begin
      RAM[RAM_MPORT_124_addr] <= RAM_MPORT_124_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_125_en & RAM_MPORT_125_mask) begin
      RAM[RAM_MPORT_125_addr] <= RAM_MPORT_125_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_126_en & RAM_MPORT_126_mask) begin
      RAM[RAM_MPORT_126_addr] <= RAM_MPORT_126_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_127_en & RAM_MPORT_127_mask) begin
      RAM[RAM_MPORT_127_addr] <= RAM_MPORT_127_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_128_en & RAM_MPORT_128_mask) begin
      RAM[RAM_MPORT_128_addr] <= RAM_MPORT_128_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_129_en & RAM_MPORT_129_mask) begin
      RAM[RAM_MPORT_129_addr] <= RAM_MPORT_129_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_130_en & RAM_MPORT_130_mask) begin
      RAM[RAM_MPORT_130_addr] <= RAM_MPORT_130_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_131_en & RAM_MPORT_131_mask) begin
      RAM[RAM_MPORT_131_addr] <= RAM_MPORT_131_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_132_en & RAM_MPORT_132_mask) begin
      RAM[RAM_MPORT_132_addr] <= RAM_MPORT_132_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_133_en & RAM_MPORT_133_mask) begin
      RAM[RAM_MPORT_133_addr] <= RAM_MPORT_133_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_134_en & RAM_MPORT_134_mask) begin
      RAM[RAM_MPORT_134_addr] <= RAM_MPORT_134_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_135_en & RAM_MPORT_135_mask) begin
      RAM[RAM_MPORT_135_addr] <= RAM_MPORT_135_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_136_en & RAM_MPORT_136_mask) begin
      RAM[RAM_MPORT_136_addr] <= RAM_MPORT_136_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_137_en & RAM_MPORT_137_mask) begin
      RAM[RAM_MPORT_137_addr] <= RAM_MPORT_137_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_138_en & RAM_MPORT_138_mask) begin
      RAM[RAM_MPORT_138_addr] <= RAM_MPORT_138_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_139_en & RAM_MPORT_139_mask) begin
      RAM[RAM_MPORT_139_addr] <= RAM_MPORT_139_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_140_en & RAM_MPORT_140_mask) begin
      RAM[RAM_MPORT_140_addr] <= RAM_MPORT_140_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_141_en & RAM_MPORT_141_mask) begin
      RAM[RAM_MPORT_141_addr] <= RAM_MPORT_141_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_142_en & RAM_MPORT_142_mask) begin
      RAM[RAM_MPORT_142_addr] <= RAM_MPORT_142_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_143_en & RAM_MPORT_143_mask) begin
      RAM[RAM_MPORT_143_addr] <= RAM_MPORT_143_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_144_en & RAM_MPORT_144_mask) begin
      RAM[RAM_MPORT_144_addr] <= RAM_MPORT_144_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_145_en & RAM_MPORT_145_mask) begin
      RAM[RAM_MPORT_145_addr] <= RAM_MPORT_145_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_146_en & RAM_MPORT_146_mask) begin
      RAM[RAM_MPORT_146_addr] <= RAM_MPORT_146_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_147_en & RAM_MPORT_147_mask) begin
      RAM[RAM_MPORT_147_addr] <= RAM_MPORT_147_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_148_en & RAM_MPORT_148_mask) begin
      RAM[RAM_MPORT_148_addr] <= RAM_MPORT_148_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_149_en & RAM_MPORT_149_mask) begin
      RAM[RAM_MPORT_149_addr] <= RAM_MPORT_149_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_150_en & RAM_MPORT_150_mask) begin
      RAM[RAM_MPORT_150_addr] <= RAM_MPORT_150_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_151_en & RAM_MPORT_151_mask) begin
      RAM[RAM_MPORT_151_addr] <= RAM_MPORT_151_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_152_en & RAM_MPORT_152_mask) begin
      RAM[RAM_MPORT_152_addr] <= RAM_MPORT_152_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_153_en & RAM_MPORT_153_mask) begin
      RAM[RAM_MPORT_153_addr] <= RAM_MPORT_153_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_154_en & RAM_MPORT_154_mask) begin
      RAM[RAM_MPORT_154_addr] <= RAM_MPORT_154_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_155_en & RAM_MPORT_155_mask) begin
      RAM[RAM_MPORT_155_addr] <= RAM_MPORT_155_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_156_en & RAM_MPORT_156_mask) begin
      RAM[RAM_MPORT_156_addr] <= RAM_MPORT_156_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_157_en & RAM_MPORT_157_mask) begin
      RAM[RAM_MPORT_157_addr] <= RAM_MPORT_157_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_158_en & RAM_MPORT_158_mask) begin
      RAM[RAM_MPORT_158_addr] <= RAM_MPORT_158_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_159_en & RAM_MPORT_159_mask) begin
      RAM[RAM_MPORT_159_addr] <= RAM_MPORT_159_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_160_en & RAM_MPORT_160_mask) begin
      RAM[RAM_MPORT_160_addr] <= RAM_MPORT_160_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_161_en & RAM_MPORT_161_mask) begin
      RAM[RAM_MPORT_161_addr] <= RAM_MPORT_161_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_162_en & RAM_MPORT_162_mask) begin
      RAM[RAM_MPORT_162_addr] <= RAM_MPORT_162_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_163_en & RAM_MPORT_163_mask) begin
      RAM[RAM_MPORT_163_addr] <= RAM_MPORT_163_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_164_en & RAM_MPORT_164_mask) begin
      RAM[RAM_MPORT_164_addr] <= RAM_MPORT_164_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_165_en & RAM_MPORT_165_mask) begin
      RAM[RAM_MPORT_165_addr] <= RAM_MPORT_165_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_166_en & RAM_MPORT_166_mask) begin
      RAM[RAM_MPORT_166_addr] <= RAM_MPORT_166_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_167_en & RAM_MPORT_167_mask) begin
      RAM[RAM_MPORT_167_addr] <= RAM_MPORT_167_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_168_en & RAM_MPORT_168_mask) begin
      RAM[RAM_MPORT_168_addr] <= RAM_MPORT_168_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_169_en & RAM_MPORT_169_mask) begin
      RAM[RAM_MPORT_169_addr] <= RAM_MPORT_169_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_170_en & RAM_MPORT_170_mask) begin
      RAM[RAM_MPORT_170_addr] <= RAM_MPORT_170_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_171_en & RAM_MPORT_171_mask) begin
      RAM[RAM_MPORT_171_addr] <= RAM_MPORT_171_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_172_en & RAM_MPORT_172_mask) begin
      RAM[RAM_MPORT_172_addr] <= RAM_MPORT_172_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_173_en & RAM_MPORT_173_mask) begin
      RAM[RAM_MPORT_173_addr] <= RAM_MPORT_173_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_174_en & RAM_MPORT_174_mask) begin
      RAM[RAM_MPORT_174_addr] <= RAM_MPORT_174_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_175_en & RAM_MPORT_175_mask) begin
      RAM[RAM_MPORT_175_addr] <= RAM_MPORT_175_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_176_en & RAM_MPORT_176_mask) begin
      RAM[RAM_MPORT_176_addr] <= RAM_MPORT_176_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_177_en & RAM_MPORT_177_mask) begin
      RAM[RAM_MPORT_177_addr] <= RAM_MPORT_177_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_178_en & RAM_MPORT_178_mask) begin
      RAM[RAM_MPORT_178_addr] <= RAM_MPORT_178_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_179_en & RAM_MPORT_179_mask) begin
      RAM[RAM_MPORT_179_addr] <= RAM_MPORT_179_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_180_en & RAM_MPORT_180_mask) begin
      RAM[RAM_MPORT_180_addr] <= RAM_MPORT_180_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_181_en & RAM_MPORT_181_mask) begin
      RAM[RAM_MPORT_181_addr] <= RAM_MPORT_181_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_182_en & RAM_MPORT_182_mask) begin
      RAM[RAM_MPORT_182_addr] <= RAM_MPORT_182_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_183_en & RAM_MPORT_183_mask) begin
      RAM[RAM_MPORT_183_addr] <= RAM_MPORT_183_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_184_en & RAM_MPORT_184_mask) begin
      RAM[RAM_MPORT_184_addr] <= RAM_MPORT_184_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_185_en & RAM_MPORT_185_mask) begin
      RAM[RAM_MPORT_185_addr] <= RAM_MPORT_185_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_186_en & RAM_MPORT_186_mask) begin
      RAM[RAM_MPORT_186_addr] <= RAM_MPORT_186_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_187_en & RAM_MPORT_187_mask) begin
      RAM[RAM_MPORT_187_addr] <= RAM_MPORT_187_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_188_en & RAM_MPORT_188_mask) begin
      RAM[RAM_MPORT_188_addr] <= RAM_MPORT_188_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_189_en & RAM_MPORT_189_mask) begin
      RAM[RAM_MPORT_189_addr] <= RAM_MPORT_189_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_190_en & RAM_MPORT_190_mask) begin
      RAM[RAM_MPORT_190_addr] <= RAM_MPORT_190_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_191_en & RAM_MPORT_191_mask) begin
      RAM[RAM_MPORT_191_addr] <= RAM_MPORT_191_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_192_en & RAM_MPORT_192_mask) begin
      RAM[RAM_MPORT_192_addr] <= RAM_MPORT_192_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_193_en & RAM_MPORT_193_mask) begin
      RAM[RAM_MPORT_193_addr] <= RAM_MPORT_193_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_194_en & RAM_MPORT_194_mask) begin
      RAM[RAM_MPORT_194_addr] <= RAM_MPORT_194_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_195_en & RAM_MPORT_195_mask) begin
      RAM[RAM_MPORT_195_addr] <= RAM_MPORT_195_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_196_en & RAM_MPORT_196_mask) begin
      RAM[RAM_MPORT_196_addr] <= RAM_MPORT_196_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_197_en & RAM_MPORT_197_mask) begin
      RAM[RAM_MPORT_197_addr] <= RAM_MPORT_197_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_198_en & RAM_MPORT_198_mask) begin
      RAM[RAM_MPORT_198_addr] <= RAM_MPORT_198_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_199_en & RAM_MPORT_199_mask) begin
      RAM[RAM_MPORT_199_addr] <= RAM_MPORT_199_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_200_en & RAM_MPORT_200_mask) begin
      RAM[RAM_MPORT_200_addr] <= RAM_MPORT_200_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_201_en & RAM_MPORT_201_mask) begin
      RAM[RAM_MPORT_201_addr] <= RAM_MPORT_201_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_202_en & RAM_MPORT_202_mask) begin
      RAM[RAM_MPORT_202_addr] <= RAM_MPORT_202_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_203_en & RAM_MPORT_203_mask) begin
      RAM[RAM_MPORT_203_addr] <= RAM_MPORT_203_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_204_en & RAM_MPORT_204_mask) begin
      RAM[RAM_MPORT_204_addr] <= RAM_MPORT_204_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_205_en & RAM_MPORT_205_mask) begin
      RAM[RAM_MPORT_205_addr] <= RAM_MPORT_205_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_206_en & RAM_MPORT_206_mask) begin
      RAM[RAM_MPORT_206_addr] <= RAM_MPORT_206_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_207_en & RAM_MPORT_207_mask) begin
      RAM[RAM_MPORT_207_addr] <= RAM_MPORT_207_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_208_en & RAM_MPORT_208_mask) begin
      RAM[RAM_MPORT_208_addr] <= RAM_MPORT_208_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_209_en & RAM_MPORT_209_mask) begin
      RAM[RAM_MPORT_209_addr] <= RAM_MPORT_209_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_210_en & RAM_MPORT_210_mask) begin
      RAM[RAM_MPORT_210_addr] <= RAM_MPORT_210_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_211_en & RAM_MPORT_211_mask) begin
      RAM[RAM_MPORT_211_addr] <= RAM_MPORT_211_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_212_en & RAM_MPORT_212_mask) begin
      RAM[RAM_MPORT_212_addr] <= RAM_MPORT_212_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_213_en & RAM_MPORT_213_mask) begin
      RAM[RAM_MPORT_213_addr] <= RAM_MPORT_213_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_214_en & RAM_MPORT_214_mask) begin
      RAM[RAM_MPORT_214_addr] <= RAM_MPORT_214_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_215_en & RAM_MPORT_215_mask) begin
      RAM[RAM_MPORT_215_addr] <= RAM_MPORT_215_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_216_en & RAM_MPORT_216_mask) begin
      RAM[RAM_MPORT_216_addr] <= RAM_MPORT_216_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_217_en & RAM_MPORT_217_mask) begin
      RAM[RAM_MPORT_217_addr] <= RAM_MPORT_217_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_218_en & RAM_MPORT_218_mask) begin
      RAM[RAM_MPORT_218_addr] <= RAM_MPORT_218_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_219_en & RAM_MPORT_219_mask) begin
      RAM[RAM_MPORT_219_addr] <= RAM_MPORT_219_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_220_en & RAM_MPORT_220_mask) begin
      RAM[RAM_MPORT_220_addr] <= RAM_MPORT_220_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_221_en & RAM_MPORT_221_mask) begin
      RAM[RAM_MPORT_221_addr] <= RAM_MPORT_221_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_222_en & RAM_MPORT_222_mask) begin
      RAM[RAM_MPORT_222_addr] <= RAM_MPORT_222_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_223_en & RAM_MPORT_223_mask) begin
      RAM[RAM_MPORT_223_addr] <= RAM_MPORT_223_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_224_en & RAM_MPORT_224_mask) begin
      RAM[RAM_MPORT_224_addr] <= RAM_MPORT_224_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_225_en & RAM_MPORT_225_mask) begin
      RAM[RAM_MPORT_225_addr] <= RAM_MPORT_225_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_226_en & RAM_MPORT_226_mask) begin
      RAM[RAM_MPORT_226_addr] <= RAM_MPORT_226_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_227_en & RAM_MPORT_227_mask) begin
      RAM[RAM_MPORT_227_addr] <= RAM_MPORT_227_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_228_en & RAM_MPORT_228_mask) begin
      RAM[RAM_MPORT_228_addr] <= RAM_MPORT_228_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_229_en & RAM_MPORT_229_mask) begin
      RAM[RAM_MPORT_229_addr] <= RAM_MPORT_229_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_230_en & RAM_MPORT_230_mask) begin
      RAM[RAM_MPORT_230_addr] <= RAM_MPORT_230_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_231_en & RAM_MPORT_231_mask) begin
      RAM[RAM_MPORT_231_addr] <= RAM_MPORT_231_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_232_en & RAM_MPORT_232_mask) begin
      RAM[RAM_MPORT_232_addr] <= RAM_MPORT_232_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_233_en & RAM_MPORT_233_mask) begin
      RAM[RAM_MPORT_233_addr] <= RAM_MPORT_233_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_234_en & RAM_MPORT_234_mask) begin
      RAM[RAM_MPORT_234_addr] <= RAM_MPORT_234_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_235_en & RAM_MPORT_235_mask) begin
      RAM[RAM_MPORT_235_addr] <= RAM_MPORT_235_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_236_en & RAM_MPORT_236_mask) begin
      RAM[RAM_MPORT_236_addr] <= RAM_MPORT_236_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_237_en & RAM_MPORT_237_mask) begin
      RAM[RAM_MPORT_237_addr] <= RAM_MPORT_237_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_238_en & RAM_MPORT_238_mask) begin
      RAM[RAM_MPORT_238_addr] <= RAM_MPORT_238_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_239_en & RAM_MPORT_239_mask) begin
      RAM[RAM_MPORT_239_addr] <= RAM_MPORT_239_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_240_en & RAM_MPORT_240_mask) begin
      RAM[RAM_MPORT_240_addr] <= RAM_MPORT_240_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_241_en & RAM_MPORT_241_mask) begin
      RAM[RAM_MPORT_241_addr] <= RAM_MPORT_241_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_242_en & RAM_MPORT_242_mask) begin
      RAM[RAM_MPORT_242_addr] <= RAM_MPORT_242_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_243_en & RAM_MPORT_243_mask) begin
      RAM[RAM_MPORT_243_addr] <= RAM_MPORT_243_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_244_en & RAM_MPORT_244_mask) begin
      RAM[RAM_MPORT_244_addr] <= RAM_MPORT_244_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_245_en & RAM_MPORT_245_mask) begin
      RAM[RAM_MPORT_245_addr] <= RAM_MPORT_245_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_246_en & RAM_MPORT_246_mask) begin
      RAM[RAM_MPORT_246_addr] <= RAM_MPORT_246_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_247_en & RAM_MPORT_247_mask) begin
      RAM[RAM_MPORT_247_addr] <= RAM_MPORT_247_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_248_en & RAM_MPORT_248_mask) begin
      RAM[RAM_MPORT_248_addr] <= RAM_MPORT_248_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_249_en & RAM_MPORT_249_mask) begin
      RAM[RAM_MPORT_249_addr] <= RAM_MPORT_249_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_250_en & RAM_MPORT_250_mask) begin
      RAM[RAM_MPORT_250_addr] <= RAM_MPORT_250_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_251_en & RAM_MPORT_251_mask) begin
      RAM[RAM_MPORT_251_addr] <= RAM_MPORT_251_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_252_en & RAM_MPORT_252_mask) begin
      RAM[RAM_MPORT_252_addr] <= RAM_MPORT_252_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_253_en & RAM_MPORT_253_mask) begin
      RAM[RAM_MPORT_253_addr] <= RAM_MPORT_253_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_254_en & RAM_MPORT_254_mask) begin
      RAM[RAM_MPORT_254_addr] <= RAM_MPORT_254_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_255_en & RAM_MPORT_255_mask) begin
      RAM[RAM_MPORT_255_addr] <= RAM_MPORT_255_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_256_en & RAM_MPORT_256_mask) begin
      RAM[RAM_MPORT_256_addr] <= RAM_MPORT_256_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_257_en & RAM_MPORT_257_mask) begin
      RAM[RAM_MPORT_257_addr] <= RAM_MPORT_257_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_258_en & RAM_MPORT_258_mask) begin
      RAM[RAM_MPORT_258_addr] <= RAM_MPORT_258_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_259_en & RAM_MPORT_259_mask) begin
      RAM[RAM_MPORT_259_addr] <= RAM_MPORT_259_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_260_en & RAM_MPORT_260_mask) begin
      RAM[RAM_MPORT_260_addr] <= RAM_MPORT_260_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_261_en & RAM_MPORT_261_mask) begin
      RAM[RAM_MPORT_261_addr] <= RAM_MPORT_261_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_262_en & RAM_MPORT_262_mask) begin
      RAM[RAM_MPORT_262_addr] <= RAM_MPORT_262_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_263_en & RAM_MPORT_263_mask) begin
      RAM[RAM_MPORT_263_addr] <= RAM_MPORT_263_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_264_en & RAM_MPORT_264_mask) begin
      RAM[RAM_MPORT_264_addr] <= RAM_MPORT_264_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_265_en & RAM_MPORT_265_mask) begin
      RAM[RAM_MPORT_265_addr] <= RAM_MPORT_265_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_266_en & RAM_MPORT_266_mask) begin
      RAM[RAM_MPORT_266_addr] <= RAM_MPORT_266_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_267_en & RAM_MPORT_267_mask) begin
      RAM[RAM_MPORT_267_addr] <= RAM_MPORT_267_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_268_en & RAM_MPORT_268_mask) begin
      RAM[RAM_MPORT_268_addr] <= RAM_MPORT_268_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_269_en & RAM_MPORT_269_mask) begin
      RAM[RAM_MPORT_269_addr] <= RAM_MPORT_269_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_270_en & RAM_MPORT_270_mask) begin
      RAM[RAM_MPORT_270_addr] <= RAM_MPORT_270_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_271_en & RAM_MPORT_271_mask) begin
      RAM[RAM_MPORT_271_addr] <= RAM_MPORT_271_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_272_en & RAM_MPORT_272_mask) begin
      RAM[RAM_MPORT_272_addr] <= RAM_MPORT_272_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_273_en & RAM_MPORT_273_mask) begin
      RAM[RAM_MPORT_273_addr] <= RAM_MPORT_273_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_274_en & RAM_MPORT_274_mask) begin
      RAM[RAM_MPORT_274_addr] <= RAM_MPORT_274_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_275_en & RAM_MPORT_275_mask) begin
      RAM[RAM_MPORT_275_addr] <= RAM_MPORT_275_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_276_en & RAM_MPORT_276_mask) begin
      RAM[RAM_MPORT_276_addr] <= RAM_MPORT_276_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_277_en & RAM_MPORT_277_mask) begin
      RAM[RAM_MPORT_277_addr] <= RAM_MPORT_277_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_278_en & RAM_MPORT_278_mask) begin
      RAM[RAM_MPORT_278_addr] <= RAM_MPORT_278_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_279_en & RAM_MPORT_279_mask) begin
      RAM[RAM_MPORT_279_addr] <= RAM_MPORT_279_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_280_en & RAM_MPORT_280_mask) begin
      RAM[RAM_MPORT_280_addr] <= RAM_MPORT_280_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_281_en & RAM_MPORT_281_mask) begin
      RAM[RAM_MPORT_281_addr] <= RAM_MPORT_281_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_282_en & RAM_MPORT_282_mask) begin
      RAM[RAM_MPORT_282_addr] <= RAM_MPORT_282_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_283_en & RAM_MPORT_283_mask) begin
      RAM[RAM_MPORT_283_addr] <= RAM_MPORT_283_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_284_en & RAM_MPORT_284_mask) begin
      RAM[RAM_MPORT_284_addr] <= RAM_MPORT_284_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_285_en & RAM_MPORT_285_mask) begin
      RAM[RAM_MPORT_285_addr] <= RAM_MPORT_285_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_286_en & RAM_MPORT_286_mask) begin
      RAM[RAM_MPORT_286_addr] <= RAM_MPORT_286_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_287_en & RAM_MPORT_287_mask) begin
      RAM[RAM_MPORT_287_addr] <= RAM_MPORT_287_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_288_en & RAM_MPORT_288_mask) begin
      RAM[RAM_MPORT_288_addr] <= RAM_MPORT_288_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_289_en & RAM_MPORT_289_mask) begin
      RAM[RAM_MPORT_289_addr] <= RAM_MPORT_289_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_290_en & RAM_MPORT_290_mask) begin
      RAM[RAM_MPORT_290_addr] <= RAM_MPORT_290_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_291_en & RAM_MPORT_291_mask) begin
      RAM[RAM_MPORT_291_addr] <= RAM_MPORT_291_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_292_en & RAM_MPORT_292_mask) begin
      RAM[RAM_MPORT_292_addr] <= RAM_MPORT_292_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_293_en & RAM_MPORT_293_mask) begin
      RAM[RAM_MPORT_293_addr] <= RAM_MPORT_293_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_294_en & RAM_MPORT_294_mask) begin
      RAM[RAM_MPORT_294_addr] <= RAM_MPORT_294_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_295_en & RAM_MPORT_295_mask) begin
      RAM[RAM_MPORT_295_addr] <= RAM_MPORT_295_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_296_en & RAM_MPORT_296_mask) begin
      RAM[RAM_MPORT_296_addr] <= RAM_MPORT_296_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_297_en & RAM_MPORT_297_mask) begin
      RAM[RAM_MPORT_297_addr] <= RAM_MPORT_297_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_298_en & RAM_MPORT_298_mask) begin
      RAM[RAM_MPORT_298_addr] <= RAM_MPORT_298_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_299_en & RAM_MPORT_299_mask) begin
      RAM[RAM_MPORT_299_addr] <= RAM_MPORT_299_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_300_en & RAM_MPORT_300_mask) begin
      RAM[RAM_MPORT_300_addr] <= RAM_MPORT_300_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_301_en & RAM_MPORT_301_mask) begin
      RAM[RAM_MPORT_301_addr] <= RAM_MPORT_301_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_302_en & RAM_MPORT_302_mask) begin
      RAM[RAM_MPORT_302_addr] <= RAM_MPORT_302_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_303_en & RAM_MPORT_303_mask) begin
      RAM[RAM_MPORT_303_addr] <= RAM_MPORT_303_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_304_en & RAM_MPORT_304_mask) begin
      RAM[RAM_MPORT_304_addr] <= RAM_MPORT_304_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_305_en & RAM_MPORT_305_mask) begin
      RAM[RAM_MPORT_305_addr] <= RAM_MPORT_305_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_306_en & RAM_MPORT_306_mask) begin
      RAM[RAM_MPORT_306_addr] <= RAM_MPORT_306_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_307_en & RAM_MPORT_307_mask) begin
      RAM[RAM_MPORT_307_addr] <= RAM_MPORT_307_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_308_en & RAM_MPORT_308_mask) begin
      RAM[RAM_MPORT_308_addr] <= RAM_MPORT_308_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_309_en & RAM_MPORT_309_mask) begin
      RAM[RAM_MPORT_309_addr] <= RAM_MPORT_309_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_310_en & RAM_MPORT_310_mask) begin
      RAM[RAM_MPORT_310_addr] <= RAM_MPORT_310_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_311_en & RAM_MPORT_311_mask) begin
      RAM[RAM_MPORT_311_addr] <= RAM_MPORT_311_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_312_en & RAM_MPORT_312_mask) begin
      RAM[RAM_MPORT_312_addr] <= RAM_MPORT_312_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_313_en & RAM_MPORT_313_mask) begin
      RAM[RAM_MPORT_313_addr] <= RAM_MPORT_313_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_314_en & RAM_MPORT_314_mask) begin
      RAM[RAM_MPORT_314_addr] <= RAM_MPORT_314_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_315_en & RAM_MPORT_315_mask) begin
      RAM[RAM_MPORT_315_addr] <= RAM_MPORT_315_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_316_en & RAM_MPORT_316_mask) begin
      RAM[RAM_MPORT_316_addr] <= RAM_MPORT_316_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_317_en & RAM_MPORT_317_mask) begin
      RAM[RAM_MPORT_317_addr] <= RAM_MPORT_317_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_318_en & RAM_MPORT_318_mask) begin
      RAM[RAM_MPORT_318_addr] <= RAM_MPORT_318_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_319_en & RAM_MPORT_319_mask) begin
      RAM[RAM_MPORT_319_addr] <= RAM_MPORT_319_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_320_en & RAM_MPORT_320_mask) begin
      RAM[RAM_MPORT_320_addr] <= RAM_MPORT_320_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_321_en & RAM_MPORT_321_mask) begin
      RAM[RAM_MPORT_321_addr] <= RAM_MPORT_321_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_322_en & RAM_MPORT_322_mask) begin
      RAM[RAM_MPORT_322_addr] <= RAM_MPORT_322_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_323_en & RAM_MPORT_323_mask) begin
      RAM[RAM_MPORT_323_addr] <= RAM_MPORT_323_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_324_en & RAM_MPORT_324_mask) begin
      RAM[RAM_MPORT_324_addr] <= RAM_MPORT_324_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_325_en & RAM_MPORT_325_mask) begin
      RAM[RAM_MPORT_325_addr] <= RAM_MPORT_325_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_326_en & RAM_MPORT_326_mask) begin
      RAM[RAM_MPORT_326_addr] <= RAM_MPORT_326_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_327_en & RAM_MPORT_327_mask) begin
      RAM[RAM_MPORT_327_addr] <= RAM_MPORT_327_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_328_en & RAM_MPORT_328_mask) begin
      RAM[RAM_MPORT_328_addr] <= RAM_MPORT_328_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_329_en & RAM_MPORT_329_mask) begin
      RAM[RAM_MPORT_329_addr] <= RAM_MPORT_329_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_330_en & RAM_MPORT_330_mask) begin
      RAM[RAM_MPORT_330_addr] <= RAM_MPORT_330_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_331_en & RAM_MPORT_331_mask) begin
      RAM[RAM_MPORT_331_addr] <= RAM_MPORT_331_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_332_en & RAM_MPORT_332_mask) begin
      RAM[RAM_MPORT_332_addr] <= RAM_MPORT_332_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_333_en & RAM_MPORT_333_mask) begin
      RAM[RAM_MPORT_333_addr] <= RAM_MPORT_333_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_334_en & RAM_MPORT_334_mask) begin
      RAM[RAM_MPORT_334_addr] <= RAM_MPORT_334_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_335_en & RAM_MPORT_335_mask) begin
      RAM[RAM_MPORT_335_addr] <= RAM_MPORT_335_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_336_en & RAM_MPORT_336_mask) begin
      RAM[RAM_MPORT_336_addr] <= RAM_MPORT_336_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_337_en & RAM_MPORT_337_mask) begin
      RAM[RAM_MPORT_337_addr] <= RAM_MPORT_337_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_338_en & RAM_MPORT_338_mask) begin
      RAM[RAM_MPORT_338_addr] <= RAM_MPORT_338_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_339_en & RAM_MPORT_339_mask) begin
      RAM[RAM_MPORT_339_addr] <= RAM_MPORT_339_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_340_en & RAM_MPORT_340_mask) begin
      RAM[RAM_MPORT_340_addr] <= RAM_MPORT_340_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_341_en & RAM_MPORT_341_mask) begin
      RAM[RAM_MPORT_341_addr] <= RAM_MPORT_341_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_342_en & RAM_MPORT_342_mask) begin
      RAM[RAM_MPORT_342_addr] <= RAM_MPORT_342_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_343_en & RAM_MPORT_343_mask) begin
      RAM[RAM_MPORT_343_addr] <= RAM_MPORT_343_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_344_en & RAM_MPORT_344_mask) begin
      RAM[RAM_MPORT_344_addr] <= RAM_MPORT_344_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_345_en & RAM_MPORT_345_mask) begin
      RAM[RAM_MPORT_345_addr] <= RAM_MPORT_345_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_346_en & RAM_MPORT_346_mask) begin
      RAM[RAM_MPORT_346_addr] <= RAM_MPORT_346_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_347_en & RAM_MPORT_347_mask) begin
      RAM[RAM_MPORT_347_addr] <= RAM_MPORT_347_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_348_en & RAM_MPORT_348_mask) begin
      RAM[RAM_MPORT_348_addr] <= RAM_MPORT_348_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_349_en & RAM_MPORT_349_mask) begin
      RAM[RAM_MPORT_349_addr] <= RAM_MPORT_349_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_350_en & RAM_MPORT_350_mask) begin
      RAM[RAM_MPORT_350_addr] <= RAM_MPORT_350_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_351_en & RAM_MPORT_351_mask) begin
      RAM[RAM_MPORT_351_addr] <= RAM_MPORT_351_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_352_en & RAM_MPORT_352_mask) begin
      RAM[RAM_MPORT_352_addr] <= RAM_MPORT_352_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_353_en & RAM_MPORT_353_mask) begin
      RAM[RAM_MPORT_353_addr] <= RAM_MPORT_353_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_354_en & RAM_MPORT_354_mask) begin
      RAM[RAM_MPORT_354_addr] <= RAM_MPORT_354_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_355_en & RAM_MPORT_355_mask) begin
      RAM[RAM_MPORT_355_addr] <= RAM_MPORT_355_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_356_en & RAM_MPORT_356_mask) begin
      RAM[RAM_MPORT_356_addr] <= RAM_MPORT_356_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_357_en & RAM_MPORT_357_mask) begin
      RAM[RAM_MPORT_357_addr] <= RAM_MPORT_357_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_358_en & RAM_MPORT_358_mask) begin
      RAM[RAM_MPORT_358_addr] <= RAM_MPORT_358_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_359_en & RAM_MPORT_359_mask) begin
      RAM[RAM_MPORT_359_addr] <= RAM_MPORT_359_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_360_en & RAM_MPORT_360_mask) begin
      RAM[RAM_MPORT_360_addr] <= RAM_MPORT_360_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_361_en & RAM_MPORT_361_mask) begin
      RAM[RAM_MPORT_361_addr] <= RAM_MPORT_361_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_362_en & RAM_MPORT_362_mask) begin
      RAM[RAM_MPORT_362_addr] <= RAM_MPORT_362_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_363_en & RAM_MPORT_363_mask) begin
      RAM[RAM_MPORT_363_addr] <= RAM_MPORT_363_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_364_en & RAM_MPORT_364_mask) begin
      RAM[RAM_MPORT_364_addr] <= RAM_MPORT_364_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_365_en & RAM_MPORT_365_mask) begin
      RAM[RAM_MPORT_365_addr] <= RAM_MPORT_365_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_366_en & RAM_MPORT_366_mask) begin
      RAM[RAM_MPORT_366_addr] <= RAM_MPORT_366_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_367_en & RAM_MPORT_367_mask) begin
      RAM[RAM_MPORT_367_addr] <= RAM_MPORT_367_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_368_en & RAM_MPORT_368_mask) begin
      RAM[RAM_MPORT_368_addr] <= RAM_MPORT_368_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_369_en & RAM_MPORT_369_mask) begin
      RAM[RAM_MPORT_369_addr] <= RAM_MPORT_369_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_370_en & RAM_MPORT_370_mask) begin
      RAM[RAM_MPORT_370_addr] <= RAM_MPORT_370_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_371_en & RAM_MPORT_371_mask) begin
      RAM[RAM_MPORT_371_addr] <= RAM_MPORT_371_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_372_en & RAM_MPORT_372_mask) begin
      RAM[RAM_MPORT_372_addr] <= RAM_MPORT_372_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_373_en & RAM_MPORT_373_mask) begin
      RAM[RAM_MPORT_373_addr] <= RAM_MPORT_373_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_374_en & RAM_MPORT_374_mask) begin
      RAM[RAM_MPORT_374_addr] <= RAM_MPORT_374_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_375_en & RAM_MPORT_375_mask) begin
      RAM[RAM_MPORT_375_addr] <= RAM_MPORT_375_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_376_en & RAM_MPORT_376_mask) begin
      RAM[RAM_MPORT_376_addr] <= RAM_MPORT_376_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_377_en & RAM_MPORT_377_mask) begin
      RAM[RAM_MPORT_377_addr] <= RAM_MPORT_377_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_378_en & RAM_MPORT_378_mask) begin
      RAM[RAM_MPORT_378_addr] <= RAM_MPORT_378_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_379_en & RAM_MPORT_379_mask) begin
      RAM[RAM_MPORT_379_addr] <= RAM_MPORT_379_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_380_en & RAM_MPORT_380_mask) begin
      RAM[RAM_MPORT_380_addr] <= RAM_MPORT_380_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_381_en & RAM_MPORT_381_mask) begin
      RAM[RAM_MPORT_381_addr] <= RAM_MPORT_381_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_382_en & RAM_MPORT_382_mask) begin
      RAM[RAM_MPORT_382_addr] <= RAM_MPORT_382_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_383_en & RAM_MPORT_383_mask) begin
      RAM[RAM_MPORT_383_addr] <= RAM_MPORT_383_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_384_en & RAM_MPORT_384_mask) begin
      RAM[RAM_MPORT_384_addr] <= RAM_MPORT_384_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_385_en & RAM_MPORT_385_mask) begin
      RAM[RAM_MPORT_385_addr] <= RAM_MPORT_385_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_386_en & RAM_MPORT_386_mask) begin
      RAM[RAM_MPORT_386_addr] <= RAM_MPORT_386_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_387_en & RAM_MPORT_387_mask) begin
      RAM[RAM_MPORT_387_addr] <= RAM_MPORT_387_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_388_en & RAM_MPORT_388_mask) begin
      RAM[RAM_MPORT_388_addr] <= RAM_MPORT_388_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_389_en & RAM_MPORT_389_mask) begin
      RAM[RAM_MPORT_389_addr] <= RAM_MPORT_389_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_390_en & RAM_MPORT_390_mask) begin
      RAM[RAM_MPORT_390_addr] <= RAM_MPORT_390_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_391_en & RAM_MPORT_391_mask) begin
      RAM[RAM_MPORT_391_addr] <= RAM_MPORT_391_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_392_en & RAM_MPORT_392_mask) begin
      RAM[RAM_MPORT_392_addr] <= RAM_MPORT_392_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_393_en & RAM_MPORT_393_mask) begin
      RAM[RAM_MPORT_393_addr] <= RAM_MPORT_393_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_394_en & RAM_MPORT_394_mask) begin
      RAM[RAM_MPORT_394_addr] <= RAM_MPORT_394_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_395_en & RAM_MPORT_395_mask) begin
      RAM[RAM_MPORT_395_addr] <= RAM_MPORT_395_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_396_en & RAM_MPORT_396_mask) begin
      RAM[RAM_MPORT_396_addr] <= RAM_MPORT_396_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_397_en & RAM_MPORT_397_mask) begin
      RAM[RAM_MPORT_397_addr] <= RAM_MPORT_397_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_398_en & RAM_MPORT_398_mask) begin
      RAM[RAM_MPORT_398_addr] <= RAM_MPORT_398_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_399_en & RAM_MPORT_399_mask) begin
      RAM[RAM_MPORT_399_addr] <= RAM_MPORT_399_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_400_en & RAM_MPORT_400_mask) begin
      RAM[RAM_MPORT_400_addr] <= RAM_MPORT_400_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_401_en & RAM_MPORT_401_mask) begin
      RAM[RAM_MPORT_401_addr] <= RAM_MPORT_401_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_402_en & RAM_MPORT_402_mask) begin
      RAM[RAM_MPORT_402_addr] <= RAM_MPORT_402_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_403_en & RAM_MPORT_403_mask) begin
      RAM[RAM_MPORT_403_addr] <= RAM_MPORT_403_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_404_en & RAM_MPORT_404_mask) begin
      RAM[RAM_MPORT_404_addr] <= RAM_MPORT_404_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_405_en & RAM_MPORT_405_mask) begin
      RAM[RAM_MPORT_405_addr] <= RAM_MPORT_405_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_406_en & RAM_MPORT_406_mask) begin
      RAM[RAM_MPORT_406_addr] <= RAM_MPORT_406_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_407_en & RAM_MPORT_407_mask) begin
      RAM[RAM_MPORT_407_addr] <= RAM_MPORT_407_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_408_en & RAM_MPORT_408_mask) begin
      RAM[RAM_MPORT_408_addr] <= RAM_MPORT_408_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_409_en & RAM_MPORT_409_mask) begin
      RAM[RAM_MPORT_409_addr] <= RAM_MPORT_409_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_410_en & RAM_MPORT_410_mask) begin
      RAM[RAM_MPORT_410_addr] <= RAM_MPORT_410_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_411_en & RAM_MPORT_411_mask) begin
      RAM[RAM_MPORT_411_addr] <= RAM_MPORT_411_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_412_en & RAM_MPORT_412_mask) begin
      RAM[RAM_MPORT_412_addr] <= RAM_MPORT_412_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_413_en & RAM_MPORT_413_mask) begin
      RAM[RAM_MPORT_413_addr] <= RAM_MPORT_413_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_414_en & RAM_MPORT_414_mask) begin
      RAM[RAM_MPORT_414_addr] <= RAM_MPORT_414_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_415_en & RAM_MPORT_415_mask) begin
      RAM[RAM_MPORT_415_addr] <= RAM_MPORT_415_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_416_en & RAM_MPORT_416_mask) begin
      RAM[RAM_MPORT_416_addr] <= RAM_MPORT_416_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_417_en & RAM_MPORT_417_mask) begin
      RAM[RAM_MPORT_417_addr] <= RAM_MPORT_417_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_418_en & RAM_MPORT_418_mask) begin
      RAM[RAM_MPORT_418_addr] <= RAM_MPORT_418_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_419_en & RAM_MPORT_419_mask) begin
      RAM[RAM_MPORT_419_addr] <= RAM_MPORT_419_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_420_en & RAM_MPORT_420_mask) begin
      RAM[RAM_MPORT_420_addr] <= RAM_MPORT_420_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_421_en & RAM_MPORT_421_mask) begin
      RAM[RAM_MPORT_421_addr] <= RAM_MPORT_421_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_422_en & RAM_MPORT_422_mask) begin
      RAM[RAM_MPORT_422_addr] <= RAM_MPORT_422_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_423_en & RAM_MPORT_423_mask) begin
      RAM[RAM_MPORT_423_addr] <= RAM_MPORT_423_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_424_en & RAM_MPORT_424_mask) begin
      RAM[RAM_MPORT_424_addr] <= RAM_MPORT_424_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_425_en & RAM_MPORT_425_mask) begin
      RAM[RAM_MPORT_425_addr] <= RAM_MPORT_425_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_426_en & RAM_MPORT_426_mask) begin
      RAM[RAM_MPORT_426_addr] <= RAM_MPORT_426_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_427_en & RAM_MPORT_427_mask) begin
      RAM[RAM_MPORT_427_addr] <= RAM_MPORT_427_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_428_en & RAM_MPORT_428_mask) begin
      RAM[RAM_MPORT_428_addr] <= RAM_MPORT_428_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_429_en & RAM_MPORT_429_mask) begin
      RAM[RAM_MPORT_429_addr] <= RAM_MPORT_429_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_430_en & RAM_MPORT_430_mask) begin
      RAM[RAM_MPORT_430_addr] <= RAM_MPORT_430_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_431_en & RAM_MPORT_431_mask) begin
      RAM[RAM_MPORT_431_addr] <= RAM_MPORT_431_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_432_en & RAM_MPORT_432_mask) begin
      RAM[RAM_MPORT_432_addr] <= RAM_MPORT_432_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_433_en & RAM_MPORT_433_mask) begin
      RAM[RAM_MPORT_433_addr] <= RAM_MPORT_433_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_434_en & RAM_MPORT_434_mask) begin
      RAM[RAM_MPORT_434_addr] <= RAM_MPORT_434_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_435_en & RAM_MPORT_435_mask) begin
      RAM[RAM_MPORT_435_addr] <= RAM_MPORT_435_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_436_en & RAM_MPORT_436_mask) begin
      RAM[RAM_MPORT_436_addr] <= RAM_MPORT_436_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_437_en & RAM_MPORT_437_mask) begin
      RAM[RAM_MPORT_437_addr] <= RAM_MPORT_437_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_438_en & RAM_MPORT_438_mask) begin
      RAM[RAM_MPORT_438_addr] <= RAM_MPORT_438_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_439_en & RAM_MPORT_439_mask) begin
      RAM[RAM_MPORT_439_addr] <= RAM_MPORT_439_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_440_en & RAM_MPORT_440_mask) begin
      RAM[RAM_MPORT_440_addr] <= RAM_MPORT_440_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_441_en & RAM_MPORT_441_mask) begin
      RAM[RAM_MPORT_441_addr] <= RAM_MPORT_441_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_442_en & RAM_MPORT_442_mask) begin
      RAM[RAM_MPORT_442_addr] <= RAM_MPORT_442_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_443_en & RAM_MPORT_443_mask) begin
      RAM[RAM_MPORT_443_addr] <= RAM_MPORT_443_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_444_en & RAM_MPORT_444_mask) begin
      RAM[RAM_MPORT_444_addr] <= RAM_MPORT_444_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_445_en & RAM_MPORT_445_mask) begin
      RAM[RAM_MPORT_445_addr] <= RAM_MPORT_445_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_446_en & RAM_MPORT_446_mask) begin
      RAM[RAM_MPORT_446_addr] <= RAM_MPORT_446_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_447_en & RAM_MPORT_447_mask) begin
      RAM[RAM_MPORT_447_addr] <= RAM_MPORT_447_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_448_en & RAM_MPORT_448_mask) begin
      RAM[RAM_MPORT_448_addr] <= RAM_MPORT_448_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_449_en & RAM_MPORT_449_mask) begin
      RAM[RAM_MPORT_449_addr] <= RAM_MPORT_449_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_450_en & RAM_MPORT_450_mask) begin
      RAM[RAM_MPORT_450_addr] <= RAM_MPORT_450_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_451_en & RAM_MPORT_451_mask) begin
      RAM[RAM_MPORT_451_addr] <= RAM_MPORT_451_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_452_en & RAM_MPORT_452_mask) begin
      RAM[RAM_MPORT_452_addr] <= RAM_MPORT_452_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_453_en & RAM_MPORT_453_mask) begin
      RAM[RAM_MPORT_453_addr] <= RAM_MPORT_453_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_454_en & RAM_MPORT_454_mask) begin
      RAM[RAM_MPORT_454_addr] <= RAM_MPORT_454_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_455_en & RAM_MPORT_455_mask) begin
      RAM[RAM_MPORT_455_addr] <= RAM_MPORT_455_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_456_en & RAM_MPORT_456_mask) begin
      RAM[RAM_MPORT_456_addr] <= RAM_MPORT_456_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_457_en & RAM_MPORT_457_mask) begin
      RAM[RAM_MPORT_457_addr] <= RAM_MPORT_457_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_458_en & RAM_MPORT_458_mask) begin
      RAM[RAM_MPORT_458_addr] <= RAM_MPORT_458_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_459_en & RAM_MPORT_459_mask) begin
      RAM[RAM_MPORT_459_addr] <= RAM_MPORT_459_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_460_en & RAM_MPORT_460_mask) begin
      RAM[RAM_MPORT_460_addr] <= RAM_MPORT_460_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_461_en & RAM_MPORT_461_mask) begin
      RAM[RAM_MPORT_461_addr] <= RAM_MPORT_461_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_462_en & RAM_MPORT_462_mask) begin
      RAM[RAM_MPORT_462_addr] <= RAM_MPORT_462_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_463_en & RAM_MPORT_463_mask) begin
      RAM[RAM_MPORT_463_addr] <= RAM_MPORT_463_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_464_en & RAM_MPORT_464_mask) begin
      RAM[RAM_MPORT_464_addr] <= RAM_MPORT_464_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_465_en & RAM_MPORT_465_mask) begin
      RAM[RAM_MPORT_465_addr] <= RAM_MPORT_465_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_466_en & RAM_MPORT_466_mask) begin
      RAM[RAM_MPORT_466_addr] <= RAM_MPORT_466_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_467_en & RAM_MPORT_467_mask) begin
      RAM[RAM_MPORT_467_addr] <= RAM_MPORT_467_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_468_en & RAM_MPORT_468_mask) begin
      RAM[RAM_MPORT_468_addr] <= RAM_MPORT_468_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_469_en & RAM_MPORT_469_mask) begin
      RAM[RAM_MPORT_469_addr] <= RAM_MPORT_469_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_470_en & RAM_MPORT_470_mask) begin
      RAM[RAM_MPORT_470_addr] <= RAM_MPORT_470_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_471_en & RAM_MPORT_471_mask) begin
      RAM[RAM_MPORT_471_addr] <= RAM_MPORT_471_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_472_en & RAM_MPORT_472_mask) begin
      RAM[RAM_MPORT_472_addr] <= RAM_MPORT_472_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_473_en & RAM_MPORT_473_mask) begin
      RAM[RAM_MPORT_473_addr] <= RAM_MPORT_473_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_474_en & RAM_MPORT_474_mask) begin
      RAM[RAM_MPORT_474_addr] <= RAM_MPORT_474_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_475_en & RAM_MPORT_475_mask) begin
      RAM[RAM_MPORT_475_addr] <= RAM_MPORT_475_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_476_en & RAM_MPORT_476_mask) begin
      RAM[RAM_MPORT_476_addr] <= RAM_MPORT_476_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_477_en & RAM_MPORT_477_mask) begin
      RAM[RAM_MPORT_477_addr] <= RAM_MPORT_477_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_478_en & RAM_MPORT_478_mask) begin
      RAM[RAM_MPORT_478_addr] <= RAM_MPORT_478_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_479_en & RAM_MPORT_479_mask) begin
      RAM[RAM_MPORT_479_addr] <= RAM_MPORT_479_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_480_en & RAM_MPORT_480_mask) begin
      RAM[RAM_MPORT_480_addr] <= RAM_MPORT_480_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_481_en & RAM_MPORT_481_mask) begin
      RAM[RAM_MPORT_481_addr] <= RAM_MPORT_481_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_482_en & RAM_MPORT_482_mask) begin
      RAM[RAM_MPORT_482_addr] <= RAM_MPORT_482_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_483_en & RAM_MPORT_483_mask) begin
      RAM[RAM_MPORT_483_addr] <= RAM_MPORT_483_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_484_en & RAM_MPORT_484_mask) begin
      RAM[RAM_MPORT_484_addr] <= RAM_MPORT_484_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_485_en & RAM_MPORT_485_mask) begin
      RAM[RAM_MPORT_485_addr] <= RAM_MPORT_485_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_486_en & RAM_MPORT_486_mask) begin
      RAM[RAM_MPORT_486_addr] <= RAM_MPORT_486_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_487_en & RAM_MPORT_487_mask) begin
      RAM[RAM_MPORT_487_addr] <= RAM_MPORT_487_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_488_en & RAM_MPORT_488_mask) begin
      RAM[RAM_MPORT_488_addr] <= RAM_MPORT_488_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_489_en & RAM_MPORT_489_mask) begin
      RAM[RAM_MPORT_489_addr] <= RAM_MPORT_489_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_490_en & RAM_MPORT_490_mask) begin
      RAM[RAM_MPORT_490_addr] <= RAM_MPORT_490_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_491_en & RAM_MPORT_491_mask) begin
      RAM[RAM_MPORT_491_addr] <= RAM_MPORT_491_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_492_en & RAM_MPORT_492_mask) begin
      RAM[RAM_MPORT_492_addr] <= RAM_MPORT_492_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_493_en & RAM_MPORT_493_mask) begin
      RAM[RAM_MPORT_493_addr] <= RAM_MPORT_493_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_494_en & RAM_MPORT_494_mask) begin
      RAM[RAM_MPORT_494_addr] <= RAM_MPORT_494_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_495_en & RAM_MPORT_495_mask) begin
      RAM[RAM_MPORT_495_addr] <= RAM_MPORT_495_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_496_en & RAM_MPORT_496_mask) begin
      RAM[RAM_MPORT_496_addr] <= RAM_MPORT_496_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_497_en & RAM_MPORT_497_mask) begin
      RAM[RAM_MPORT_497_addr] <= RAM_MPORT_497_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_498_en & RAM_MPORT_498_mask) begin
      RAM[RAM_MPORT_498_addr] <= RAM_MPORT_498_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_499_en & RAM_MPORT_499_mask) begin
      RAM[RAM_MPORT_499_addr] <= RAM_MPORT_499_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_500_en & RAM_MPORT_500_mask) begin
      RAM[RAM_MPORT_500_addr] <= RAM_MPORT_500_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_501_en & RAM_MPORT_501_mask) begin
      RAM[RAM_MPORT_501_addr] <= RAM_MPORT_501_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_502_en & RAM_MPORT_502_mask) begin
      RAM[RAM_MPORT_502_addr] <= RAM_MPORT_502_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_503_en & RAM_MPORT_503_mask) begin
      RAM[RAM_MPORT_503_addr] <= RAM_MPORT_503_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_504_en & RAM_MPORT_504_mask) begin
      RAM[RAM_MPORT_504_addr] <= RAM_MPORT_504_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_505_en & RAM_MPORT_505_mask) begin
      RAM[RAM_MPORT_505_addr] <= RAM_MPORT_505_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_506_en & RAM_MPORT_506_mask) begin
      RAM[RAM_MPORT_506_addr] <= RAM_MPORT_506_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_507_en & RAM_MPORT_507_mask) begin
      RAM[RAM_MPORT_507_addr] <= RAM_MPORT_507_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_508_en & RAM_MPORT_508_mask) begin
      RAM[RAM_MPORT_508_addr] <= RAM_MPORT_508_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_509_en & RAM_MPORT_509_mask) begin
      RAM[RAM_MPORT_509_addr] <= RAM_MPORT_509_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_510_en & RAM_MPORT_510_mask) begin
      RAM[RAM_MPORT_510_addr] <= RAM_MPORT_510_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_511_en & RAM_MPORT_511_mask) begin
      RAM[RAM_MPORT_511_addr] <= RAM_MPORT_511_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_512_en & RAM_MPORT_512_mask) begin
      RAM[RAM_MPORT_512_addr] <= RAM_MPORT_512_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_513_en & RAM_MPORT_513_mask) begin
      RAM[RAM_MPORT_513_addr] <= RAM_MPORT_513_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_514_en & RAM_MPORT_514_mask) begin
      RAM[RAM_MPORT_514_addr] <= RAM_MPORT_514_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_515_en & RAM_MPORT_515_mask) begin
      RAM[RAM_MPORT_515_addr] <= RAM_MPORT_515_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_516_en & RAM_MPORT_516_mask) begin
      RAM[RAM_MPORT_516_addr] <= RAM_MPORT_516_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_517_en & RAM_MPORT_517_mask) begin
      RAM[RAM_MPORT_517_addr] <= RAM_MPORT_517_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_518_en & RAM_MPORT_518_mask) begin
      RAM[RAM_MPORT_518_addr] <= RAM_MPORT_518_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_519_en & RAM_MPORT_519_mask) begin
      RAM[RAM_MPORT_519_addr] <= RAM_MPORT_519_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_520_en & RAM_MPORT_520_mask) begin
      RAM[RAM_MPORT_520_addr] <= RAM_MPORT_520_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_521_en & RAM_MPORT_521_mask) begin
      RAM[RAM_MPORT_521_addr] <= RAM_MPORT_521_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_522_en & RAM_MPORT_522_mask) begin
      RAM[RAM_MPORT_522_addr] <= RAM_MPORT_522_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_523_en & RAM_MPORT_523_mask) begin
      RAM[RAM_MPORT_523_addr] <= RAM_MPORT_523_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_524_en & RAM_MPORT_524_mask) begin
      RAM[RAM_MPORT_524_addr] <= RAM_MPORT_524_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_525_en & RAM_MPORT_525_mask) begin
      RAM[RAM_MPORT_525_addr] <= RAM_MPORT_525_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_526_en & RAM_MPORT_526_mask) begin
      RAM[RAM_MPORT_526_addr] <= RAM_MPORT_526_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_527_en & RAM_MPORT_527_mask) begin
      RAM[RAM_MPORT_527_addr] <= RAM_MPORT_527_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_528_en & RAM_MPORT_528_mask) begin
      RAM[RAM_MPORT_528_addr] <= RAM_MPORT_528_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_529_en & RAM_MPORT_529_mask) begin
      RAM[RAM_MPORT_529_addr] <= RAM_MPORT_529_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_530_en & RAM_MPORT_530_mask) begin
      RAM[RAM_MPORT_530_addr] <= RAM_MPORT_530_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_531_en & RAM_MPORT_531_mask) begin
      RAM[RAM_MPORT_531_addr] <= RAM_MPORT_531_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_532_en & RAM_MPORT_532_mask) begin
      RAM[RAM_MPORT_532_addr] <= RAM_MPORT_532_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_533_en & RAM_MPORT_533_mask) begin
      RAM[RAM_MPORT_533_addr] <= RAM_MPORT_533_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_534_en & RAM_MPORT_534_mask) begin
      RAM[RAM_MPORT_534_addr] <= RAM_MPORT_534_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_535_en & RAM_MPORT_535_mask) begin
      RAM[RAM_MPORT_535_addr] <= RAM_MPORT_535_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_536_en & RAM_MPORT_536_mask) begin
      RAM[RAM_MPORT_536_addr] <= RAM_MPORT_536_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_537_en & RAM_MPORT_537_mask) begin
      RAM[RAM_MPORT_537_addr] <= RAM_MPORT_537_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_538_en & RAM_MPORT_538_mask) begin
      RAM[RAM_MPORT_538_addr] <= RAM_MPORT_538_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_539_en & RAM_MPORT_539_mask) begin
      RAM[RAM_MPORT_539_addr] <= RAM_MPORT_539_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_540_en & RAM_MPORT_540_mask) begin
      RAM[RAM_MPORT_540_addr] <= RAM_MPORT_540_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_541_en & RAM_MPORT_541_mask) begin
      RAM[RAM_MPORT_541_addr] <= RAM_MPORT_541_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_542_en & RAM_MPORT_542_mask) begin
      RAM[RAM_MPORT_542_addr] <= RAM_MPORT_542_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_543_en & RAM_MPORT_543_mask) begin
      RAM[RAM_MPORT_543_addr] <= RAM_MPORT_543_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_544_en & RAM_MPORT_544_mask) begin
      RAM[RAM_MPORT_544_addr] <= RAM_MPORT_544_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_545_en & RAM_MPORT_545_mask) begin
      RAM[RAM_MPORT_545_addr] <= RAM_MPORT_545_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_546_en & RAM_MPORT_546_mask) begin
      RAM[RAM_MPORT_546_addr] <= RAM_MPORT_546_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_547_en & RAM_MPORT_547_mask) begin
      RAM[RAM_MPORT_547_addr] <= RAM_MPORT_547_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_548_en & RAM_MPORT_548_mask) begin
      RAM[RAM_MPORT_548_addr] <= RAM_MPORT_548_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_549_en & RAM_MPORT_549_mask) begin
      RAM[RAM_MPORT_549_addr] <= RAM_MPORT_549_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_550_en & RAM_MPORT_550_mask) begin
      RAM[RAM_MPORT_550_addr] <= RAM_MPORT_550_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_551_en & RAM_MPORT_551_mask) begin
      RAM[RAM_MPORT_551_addr] <= RAM_MPORT_551_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_552_en & RAM_MPORT_552_mask) begin
      RAM[RAM_MPORT_552_addr] <= RAM_MPORT_552_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_553_en & RAM_MPORT_553_mask) begin
      RAM[RAM_MPORT_553_addr] <= RAM_MPORT_553_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_554_en & RAM_MPORT_554_mask) begin
      RAM[RAM_MPORT_554_addr] <= RAM_MPORT_554_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_555_en & RAM_MPORT_555_mask) begin
      RAM[RAM_MPORT_555_addr] <= RAM_MPORT_555_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_556_en & RAM_MPORT_556_mask) begin
      RAM[RAM_MPORT_556_addr] <= RAM_MPORT_556_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_557_en & RAM_MPORT_557_mask) begin
      RAM[RAM_MPORT_557_addr] <= RAM_MPORT_557_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_558_en & RAM_MPORT_558_mask) begin
      RAM[RAM_MPORT_558_addr] <= RAM_MPORT_558_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_559_en & RAM_MPORT_559_mask) begin
      RAM[RAM_MPORT_559_addr] <= RAM_MPORT_559_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_560_en & RAM_MPORT_560_mask) begin
      RAM[RAM_MPORT_560_addr] <= RAM_MPORT_560_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_561_en & RAM_MPORT_561_mask) begin
      RAM[RAM_MPORT_561_addr] <= RAM_MPORT_561_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_562_en & RAM_MPORT_562_mask) begin
      RAM[RAM_MPORT_562_addr] <= RAM_MPORT_562_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_563_en & RAM_MPORT_563_mask) begin
      RAM[RAM_MPORT_563_addr] <= RAM_MPORT_563_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_564_en & RAM_MPORT_564_mask) begin
      RAM[RAM_MPORT_564_addr] <= RAM_MPORT_564_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_565_en & RAM_MPORT_565_mask) begin
      RAM[RAM_MPORT_565_addr] <= RAM_MPORT_565_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_566_en & RAM_MPORT_566_mask) begin
      RAM[RAM_MPORT_566_addr] <= RAM_MPORT_566_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_567_en & RAM_MPORT_567_mask) begin
      RAM[RAM_MPORT_567_addr] <= RAM_MPORT_567_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_568_en & RAM_MPORT_568_mask) begin
      RAM[RAM_MPORT_568_addr] <= RAM_MPORT_568_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_569_en & RAM_MPORT_569_mask) begin
      RAM[RAM_MPORT_569_addr] <= RAM_MPORT_569_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_570_en & RAM_MPORT_570_mask) begin
      RAM[RAM_MPORT_570_addr] <= RAM_MPORT_570_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_571_en & RAM_MPORT_571_mask) begin
      RAM[RAM_MPORT_571_addr] <= RAM_MPORT_571_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_572_en & RAM_MPORT_572_mask) begin
      RAM[RAM_MPORT_572_addr] <= RAM_MPORT_572_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_573_en & RAM_MPORT_573_mask) begin
      RAM[RAM_MPORT_573_addr] <= RAM_MPORT_573_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_574_en & RAM_MPORT_574_mask) begin
      RAM[RAM_MPORT_574_addr] <= RAM_MPORT_574_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_575_en & RAM_MPORT_575_mask) begin
      RAM[RAM_MPORT_575_addr] <= RAM_MPORT_575_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_576_en & RAM_MPORT_576_mask) begin
      RAM[RAM_MPORT_576_addr] <= RAM_MPORT_576_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_577_en & RAM_MPORT_577_mask) begin
      RAM[RAM_MPORT_577_addr] <= RAM_MPORT_577_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_578_en & RAM_MPORT_578_mask) begin
      RAM[RAM_MPORT_578_addr] <= RAM_MPORT_578_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_579_en & RAM_MPORT_579_mask) begin
      RAM[RAM_MPORT_579_addr] <= RAM_MPORT_579_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_580_en & RAM_MPORT_580_mask) begin
      RAM[RAM_MPORT_580_addr] <= RAM_MPORT_580_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_581_en & RAM_MPORT_581_mask) begin
      RAM[RAM_MPORT_581_addr] <= RAM_MPORT_581_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_582_en & RAM_MPORT_582_mask) begin
      RAM[RAM_MPORT_582_addr] <= RAM_MPORT_582_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_583_en & RAM_MPORT_583_mask) begin
      RAM[RAM_MPORT_583_addr] <= RAM_MPORT_583_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_584_en & RAM_MPORT_584_mask) begin
      RAM[RAM_MPORT_584_addr] <= RAM_MPORT_584_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_585_en & RAM_MPORT_585_mask) begin
      RAM[RAM_MPORT_585_addr] <= RAM_MPORT_585_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_586_en & RAM_MPORT_586_mask) begin
      RAM[RAM_MPORT_586_addr] <= RAM_MPORT_586_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_587_en & RAM_MPORT_587_mask) begin
      RAM[RAM_MPORT_587_addr] <= RAM_MPORT_587_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_588_en & RAM_MPORT_588_mask) begin
      RAM[RAM_MPORT_588_addr] <= RAM_MPORT_588_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_589_en & RAM_MPORT_589_mask) begin
      RAM[RAM_MPORT_589_addr] <= RAM_MPORT_589_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_590_en & RAM_MPORT_590_mask) begin
      RAM[RAM_MPORT_590_addr] <= RAM_MPORT_590_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_591_en & RAM_MPORT_591_mask) begin
      RAM[RAM_MPORT_591_addr] <= RAM_MPORT_591_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_592_en & RAM_MPORT_592_mask) begin
      RAM[RAM_MPORT_592_addr] <= RAM_MPORT_592_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_593_en & RAM_MPORT_593_mask) begin
      RAM[RAM_MPORT_593_addr] <= RAM_MPORT_593_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_594_en & RAM_MPORT_594_mask) begin
      RAM[RAM_MPORT_594_addr] <= RAM_MPORT_594_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_595_en & RAM_MPORT_595_mask) begin
      RAM[RAM_MPORT_595_addr] <= RAM_MPORT_595_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_596_en & RAM_MPORT_596_mask) begin
      RAM[RAM_MPORT_596_addr] <= RAM_MPORT_596_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_597_en & RAM_MPORT_597_mask) begin
      RAM[RAM_MPORT_597_addr] <= RAM_MPORT_597_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_598_en & RAM_MPORT_598_mask) begin
      RAM[RAM_MPORT_598_addr] <= RAM_MPORT_598_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_599_en & RAM_MPORT_599_mask) begin
      RAM[RAM_MPORT_599_addr] <= RAM_MPORT_599_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_600_en & RAM_MPORT_600_mask) begin
      RAM[RAM_MPORT_600_addr] <= RAM_MPORT_600_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_601_en & RAM_MPORT_601_mask) begin
      RAM[RAM_MPORT_601_addr] <= RAM_MPORT_601_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_602_en & RAM_MPORT_602_mask) begin
      RAM[RAM_MPORT_602_addr] <= RAM_MPORT_602_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_603_en & RAM_MPORT_603_mask) begin
      RAM[RAM_MPORT_603_addr] <= RAM_MPORT_603_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_604_en & RAM_MPORT_604_mask) begin
      RAM[RAM_MPORT_604_addr] <= RAM_MPORT_604_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_605_en & RAM_MPORT_605_mask) begin
      RAM[RAM_MPORT_605_addr] <= RAM_MPORT_605_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_606_en & RAM_MPORT_606_mask) begin
      RAM[RAM_MPORT_606_addr] <= RAM_MPORT_606_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_607_en & RAM_MPORT_607_mask) begin
      RAM[RAM_MPORT_607_addr] <= RAM_MPORT_607_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_608_en & RAM_MPORT_608_mask) begin
      RAM[RAM_MPORT_608_addr] <= RAM_MPORT_608_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_609_en & RAM_MPORT_609_mask) begin
      RAM[RAM_MPORT_609_addr] <= RAM_MPORT_609_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_610_en & RAM_MPORT_610_mask) begin
      RAM[RAM_MPORT_610_addr] <= RAM_MPORT_610_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_611_en & RAM_MPORT_611_mask) begin
      RAM[RAM_MPORT_611_addr] <= RAM_MPORT_611_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_612_en & RAM_MPORT_612_mask) begin
      RAM[RAM_MPORT_612_addr] <= RAM_MPORT_612_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_613_en & RAM_MPORT_613_mask) begin
      RAM[RAM_MPORT_613_addr] <= RAM_MPORT_613_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_614_en & RAM_MPORT_614_mask) begin
      RAM[RAM_MPORT_614_addr] <= RAM_MPORT_614_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_615_en & RAM_MPORT_615_mask) begin
      RAM[RAM_MPORT_615_addr] <= RAM_MPORT_615_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_616_en & RAM_MPORT_616_mask) begin
      RAM[RAM_MPORT_616_addr] <= RAM_MPORT_616_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_617_en & RAM_MPORT_617_mask) begin
      RAM[RAM_MPORT_617_addr] <= RAM_MPORT_617_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_618_en & RAM_MPORT_618_mask) begin
      RAM[RAM_MPORT_618_addr] <= RAM_MPORT_618_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_619_en & RAM_MPORT_619_mask) begin
      RAM[RAM_MPORT_619_addr] <= RAM_MPORT_619_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_620_en & RAM_MPORT_620_mask) begin
      RAM[RAM_MPORT_620_addr] <= RAM_MPORT_620_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_621_en & RAM_MPORT_621_mask) begin
      RAM[RAM_MPORT_621_addr] <= RAM_MPORT_621_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_622_en & RAM_MPORT_622_mask) begin
      RAM[RAM_MPORT_622_addr] <= RAM_MPORT_622_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_623_en & RAM_MPORT_623_mask) begin
      RAM[RAM_MPORT_623_addr] <= RAM_MPORT_623_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_624_en & RAM_MPORT_624_mask) begin
      RAM[RAM_MPORT_624_addr] <= RAM_MPORT_624_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_625_en & RAM_MPORT_625_mask) begin
      RAM[RAM_MPORT_625_addr] <= RAM_MPORT_625_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_626_en & RAM_MPORT_626_mask) begin
      RAM[RAM_MPORT_626_addr] <= RAM_MPORT_626_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_627_en & RAM_MPORT_627_mask) begin
      RAM[RAM_MPORT_627_addr] <= RAM_MPORT_627_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_628_en & RAM_MPORT_628_mask) begin
      RAM[RAM_MPORT_628_addr] <= RAM_MPORT_628_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_629_en & RAM_MPORT_629_mask) begin
      RAM[RAM_MPORT_629_addr] <= RAM_MPORT_629_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_630_en & RAM_MPORT_630_mask) begin
      RAM[RAM_MPORT_630_addr] <= RAM_MPORT_630_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_631_en & RAM_MPORT_631_mask) begin
      RAM[RAM_MPORT_631_addr] <= RAM_MPORT_631_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_632_en & RAM_MPORT_632_mask) begin
      RAM[RAM_MPORT_632_addr] <= RAM_MPORT_632_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_633_en & RAM_MPORT_633_mask) begin
      RAM[RAM_MPORT_633_addr] <= RAM_MPORT_633_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_634_en & RAM_MPORT_634_mask) begin
      RAM[RAM_MPORT_634_addr] <= RAM_MPORT_634_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_635_en & RAM_MPORT_635_mask) begin
      RAM[RAM_MPORT_635_addr] <= RAM_MPORT_635_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_636_en & RAM_MPORT_636_mask) begin
      RAM[RAM_MPORT_636_addr] <= RAM_MPORT_636_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_637_en & RAM_MPORT_637_mask) begin
      RAM[RAM_MPORT_637_addr] <= RAM_MPORT_637_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_638_en & RAM_MPORT_638_mask) begin
      RAM[RAM_MPORT_638_addr] <= RAM_MPORT_638_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_639_en & RAM_MPORT_639_mask) begin
      RAM[RAM_MPORT_639_addr] <= RAM_MPORT_639_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_640_en & RAM_MPORT_640_mask) begin
      RAM[RAM_MPORT_640_addr] <= RAM_MPORT_640_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_641_en & RAM_MPORT_641_mask) begin
      RAM[RAM_MPORT_641_addr] <= RAM_MPORT_641_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_642_en & RAM_MPORT_642_mask) begin
      RAM[RAM_MPORT_642_addr] <= RAM_MPORT_642_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_643_en & RAM_MPORT_643_mask) begin
      RAM[RAM_MPORT_643_addr] <= RAM_MPORT_643_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_644_en & RAM_MPORT_644_mask) begin
      RAM[RAM_MPORT_644_addr] <= RAM_MPORT_644_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_645_en & RAM_MPORT_645_mask) begin
      RAM[RAM_MPORT_645_addr] <= RAM_MPORT_645_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_646_en & RAM_MPORT_646_mask) begin
      RAM[RAM_MPORT_646_addr] <= RAM_MPORT_646_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_647_en & RAM_MPORT_647_mask) begin
      RAM[RAM_MPORT_647_addr] <= RAM_MPORT_647_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_648_en & RAM_MPORT_648_mask) begin
      RAM[RAM_MPORT_648_addr] <= RAM_MPORT_648_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_649_en & RAM_MPORT_649_mask) begin
      RAM[RAM_MPORT_649_addr] <= RAM_MPORT_649_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_650_en & RAM_MPORT_650_mask) begin
      RAM[RAM_MPORT_650_addr] <= RAM_MPORT_650_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_651_en & RAM_MPORT_651_mask) begin
      RAM[RAM_MPORT_651_addr] <= RAM_MPORT_651_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_652_en & RAM_MPORT_652_mask) begin
      RAM[RAM_MPORT_652_addr] <= RAM_MPORT_652_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_653_en & RAM_MPORT_653_mask) begin
      RAM[RAM_MPORT_653_addr] <= RAM_MPORT_653_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_654_en & RAM_MPORT_654_mask) begin
      RAM[RAM_MPORT_654_addr] <= RAM_MPORT_654_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_655_en & RAM_MPORT_655_mask) begin
      RAM[RAM_MPORT_655_addr] <= RAM_MPORT_655_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_656_en & RAM_MPORT_656_mask) begin
      RAM[RAM_MPORT_656_addr] <= RAM_MPORT_656_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_657_en & RAM_MPORT_657_mask) begin
      RAM[RAM_MPORT_657_addr] <= RAM_MPORT_657_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_658_en & RAM_MPORT_658_mask) begin
      RAM[RAM_MPORT_658_addr] <= RAM_MPORT_658_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_659_en & RAM_MPORT_659_mask) begin
      RAM[RAM_MPORT_659_addr] <= RAM_MPORT_659_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_660_en & RAM_MPORT_660_mask) begin
      RAM[RAM_MPORT_660_addr] <= RAM_MPORT_660_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_661_en & RAM_MPORT_661_mask) begin
      RAM[RAM_MPORT_661_addr] <= RAM_MPORT_661_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_662_en & RAM_MPORT_662_mask) begin
      RAM[RAM_MPORT_662_addr] <= RAM_MPORT_662_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_663_en & RAM_MPORT_663_mask) begin
      RAM[RAM_MPORT_663_addr] <= RAM_MPORT_663_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_664_en & RAM_MPORT_664_mask) begin
      RAM[RAM_MPORT_664_addr] <= RAM_MPORT_664_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_665_en & RAM_MPORT_665_mask) begin
      RAM[RAM_MPORT_665_addr] <= RAM_MPORT_665_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_666_en & RAM_MPORT_666_mask) begin
      RAM[RAM_MPORT_666_addr] <= RAM_MPORT_666_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_667_en & RAM_MPORT_667_mask) begin
      RAM[RAM_MPORT_667_addr] <= RAM_MPORT_667_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_668_en & RAM_MPORT_668_mask) begin
      RAM[RAM_MPORT_668_addr] <= RAM_MPORT_668_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_669_en & RAM_MPORT_669_mask) begin
      RAM[RAM_MPORT_669_addr] <= RAM_MPORT_669_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_670_en & RAM_MPORT_670_mask) begin
      RAM[RAM_MPORT_670_addr] <= RAM_MPORT_670_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_671_en & RAM_MPORT_671_mask) begin
      RAM[RAM_MPORT_671_addr] <= RAM_MPORT_671_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_672_en & RAM_MPORT_672_mask) begin
      RAM[RAM_MPORT_672_addr] <= RAM_MPORT_672_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_673_en & RAM_MPORT_673_mask) begin
      RAM[RAM_MPORT_673_addr] <= RAM_MPORT_673_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_674_en & RAM_MPORT_674_mask) begin
      RAM[RAM_MPORT_674_addr] <= RAM_MPORT_674_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_675_en & RAM_MPORT_675_mask) begin
      RAM[RAM_MPORT_675_addr] <= RAM_MPORT_675_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_676_en & RAM_MPORT_676_mask) begin
      RAM[RAM_MPORT_676_addr] <= RAM_MPORT_676_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_677_en & RAM_MPORT_677_mask) begin
      RAM[RAM_MPORT_677_addr] <= RAM_MPORT_677_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_678_en & RAM_MPORT_678_mask) begin
      RAM[RAM_MPORT_678_addr] <= RAM_MPORT_678_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_679_en & RAM_MPORT_679_mask) begin
      RAM[RAM_MPORT_679_addr] <= RAM_MPORT_679_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_680_en & RAM_MPORT_680_mask) begin
      RAM[RAM_MPORT_680_addr] <= RAM_MPORT_680_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_681_en & RAM_MPORT_681_mask) begin
      RAM[RAM_MPORT_681_addr] <= RAM_MPORT_681_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_682_en & RAM_MPORT_682_mask) begin
      RAM[RAM_MPORT_682_addr] <= RAM_MPORT_682_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_683_en & RAM_MPORT_683_mask) begin
      RAM[RAM_MPORT_683_addr] <= RAM_MPORT_683_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_684_en & RAM_MPORT_684_mask) begin
      RAM[RAM_MPORT_684_addr] <= RAM_MPORT_684_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_685_en & RAM_MPORT_685_mask) begin
      RAM[RAM_MPORT_685_addr] <= RAM_MPORT_685_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_686_en & RAM_MPORT_686_mask) begin
      RAM[RAM_MPORT_686_addr] <= RAM_MPORT_686_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_687_en & RAM_MPORT_687_mask) begin
      RAM[RAM_MPORT_687_addr] <= RAM_MPORT_687_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_688_en & RAM_MPORT_688_mask) begin
      RAM[RAM_MPORT_688_addr] <= RAM_MPORT_688_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_689_en & RAM_MPORT_689_mask) begin
      RAM[RAM_MPORT_689_addr] <= RAM_MPORT_689_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_690_en & RAM_MPORT_690_mask) begin
      RAM[RAM_MPORT_690_addr] <= RAM_MPORT_690_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_691_en & RAM_MPORT_691_mask) begin
      RAM[RAM_MPORT_691_addr] <= RAM_MPORT_691_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_692_en & RAM_MPORT_692_mask) begin
      RAM[RAM_MPORT_692_addr] <= RAM_MPORT_692_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_693_en & RAM_MPORT_693_mask) begin
      RAM[RAM_MPORT_693_addr] <= RAM_MPORT_693_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_694_en & RAM_MPORT_694_mask) begin
      RAM[RAM_MPORT_694_addr] <= RAM_MPORT_694_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_695_en & RAM_MPORT_695_mask) begin
      RAM[RAM_MPORT_695_addr] <= RAM_MPORT_695_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_696_en & RAM_MPORT_696_mask) begin
      RAM[RAM_MPORT_696_addr] <= RAM_MPORT_696_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_697_en & RAM_MPORT_697_mask) begin
      RAM[RAM_MPORT_697_addr] <= RAM_MPORT_697_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_698_en & RAM_MPORT_698_mask) begin
      RAM[RAM_MPORT_698_addr] <= RAM_MPORT_698_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_699_en & RAM_MPORT_699_mask) begin
      RAM[RAM_MPORT_699_addr] <= RAM_MPORT_699_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_700_en & RAM_MPORT_700_mask) begin
      RAM[RAM_MPORT_700_addr] <= RAM_MPORT_700_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_701_en & RAM_MPORT_701_mask) begin
      RAM[RAM_MPORT_701_addr] <= RAM_MPORT_701_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_702_en & RAM_MPORT_702_mask) begin
      RAM[RAM_MPORT_702_addr] <= RAM_MPORT_702_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_703_en & RAM_MPORT_703_mask) begin
      RAM[RAM_MPORT_703_addr] <= RAM_MPORT_703_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_704_en & RAM_MPORT_704_mask) begin
      RAM[RAM_MPORT_704_addr] <= RAM_MPORT_704_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_705_en & RAM_MPORT_705_mask) begin
      RAM[RAM_MPORT_705_addr] <= RAM_MPORT_705_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_706_en & RAM_MPORT_706_mask) begin
      RAM[RAM_MPORT_706_addr] <= RAM_MPORT_706_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_707_en & RAM_MPORT_707_mask) begin
      RAM[RAM_MPORT_707_addr] <= RAM_MPORT_707_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_708_en & RAM_MPORT_708_mask) begin
      RAM[RAM_MPORT_708_addr] <= RAM_MPORT_708_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_709_en & RAM_MPORT_709_mask) begin
      RAM[RAM_MPORT_709_addr] <= RAM_MPORT_709_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_710_en & RAM_MPORT_710_mask) begin
      RAM[RAM_MPORT_710_addr] <= RAM_MPORT_710_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_711_en & RAM_MPORT_711_mask) begin
      RAM[RAM_MPORT_711_addr] <= RAM_MPORT_711_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_712_en & RAM_MPORT_712_mask) begin
      RAM[RAM_MPORT_712_addr] <= RAM_MPORT_712_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_713_en & RAM_MPORT_713_mask) begin
      RAM[RAM_MPORT_713_addr] <= RAM_MPORT_713_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_714_en & RAM_MPORT_714_mask) begin
      RAM[RAM_MPORT_714_addr] <= RAM_MPORT_714_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_715_en & RAM_MPORT_715_mask) begin
      RAM[RAM_MPORT_715_addr] <= RAM_MPORT_715_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_716_en & RAM_MPORT_716_mask) begin
      RAM[RAM_MPORT_716_addr] <= RAM_MPORT_716_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_717_en & RAM_MPORT_717_mask) begin
      RAM[RAM_MPORT_717_addr] <= RAM_MPORT_717_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_718_en & RAM_MPORT_718_mask) begin
      RAM[RAM_MPORT_718_addr] <= RAM_MPORT_718_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_719_en & RAM_MPORT_719_mask) begin
      RAM[RAM_MPORT_719_addr] <= RAM_MPORT_719_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_720_en & RAM_MPORT_720_mask) begin
      RAM[RAM_MPORT_720_addr] <= RAM_MPORT_720_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_721_en & RAM_MPORT_721_mask) begin
      RAM[RAM_MPORT_721_addr] <= RAM_MPORT_721_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_722_en & RAM_MPORT_722_mask) begin
      RAM[RAM_MPORT_722_addr] <= RAM_MPORT_722_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_723_en & RAM_MPORT_723_mask) begin
      RAM[RAM_MPORT_723_addr] <= RAM_MPORT_723_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_724_en & RAM_MPORT_724_mask) begin
      RAM[RAM_MPORT_724_addr] <= RAM_MPORT_724_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_725_en & RAM_MPORT_725_mask) begin
      RAM[RAM_MPORT_725_addr] <= RAM_MPORT_725_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_726_en & RAM_MPORT_726_mask) begin
      RAM[RAM_MPORT_726_addr] <= RAM_MPORT_726_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_727_en & RAM_MPORT_727_mask) begin
      RAM[RAM_MPORT_727_addr] <= RAM_MPORT_727_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_728_en & RAM_MPORT_728_mask) begin
      RAM[RAM_MPORT_728_addr] <= RAM_MPORT_728_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_729_en & RAM_MPORT_729_mask) begin
      RAM[RAM_MPORT_729_addr] <= RAM_MPORT_729_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_730_en & RAM_MPORT_730_mask) begin
      RAM[RAM_MPORT_730_addr] <= RAM_MPORT_730_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_731_en & RAM_MPORT_731_mask) begin
      RAM[RAM_MPORT_731_addr] <= RAM_MPORT_731_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_732_en & RAM_MPORT_732_mask) begin
      RAM[RAM_MPORT_732_addr] <= RAM_MPORT_732_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_733_en & RAM_MPORT_733_mask) begin
      RAM[RAM_MPORT_733_addr] <= RAM_MPORT_733_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_734_en & RAM_MPORT_734_mask) begin
      RAM[RAM_MPORT_734_addr] <= RAM_MPORT_734_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_735_en & RAM_MPORT_735_mask) begin
      RAM[RAM_MPORT_735_addr] <= RAM_MPORT_735_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_736_en & RAM_MPORT_736_mask) begin
      RAM[RAM_MPORT_736_addr] <= RAM_MPORT_736_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_737_en & RAM_MPORT_737_mask) begin
      RAM[RAM_MPORT_737_addr] <= RAM_MPORT_737_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_738_en & RAM_MPORT_738_mask) begin
      RAM[RAM_MPORT_738_addr] <= RAM_MPORT_738_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_739_en & RAM_MPORT_739_mask) begin
      RAM[RAM_MPORT_739_addr] <= RAM_MPORT_739_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_740_en & RAM_MPORT_740_mask) begin
      RAM[RAM_MPORT_740_addr] <= RAM_MPORT_740_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_741_en & RAM_MPORT_741_mask) begin
      RAM[RAM_MPORT_741_addr] <= RAM_MPORT_741_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_742_en & RAM_MPORT_742_mask) begin
      RAM[RAM_MPORT_742_addr] <= RAM_MPORT_742_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_743_en & RAM_MPORT_743_mask) begin
      RAM[RAM_MPORT_743_addr] <= RAM_MPORT_743_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_744_en & RAM_MPORT_744_mask) begin
      RAM[RAM_MPORT_744_addr] <= RAM_MPORT_744_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_745_en & RAM_MPORT_745_mask) begin
      RAM[RAM_MPORT_745_addr] <= RAM_MPORT_745_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_746_en & RAM_MPORT_746_mask) begin
      RAM[RAM_MPORT_746_addr] <= RAM_MPORT_746_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_747_en & RAM_MPORT_747_mask) begin
      RAM[RAM_MPORT_747_addr] <= RAM_MPORT_747_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_748_en & RAM_MPORT_748_mask) begin
      RAM[RAM_MPORT_748_addr] <= RAM_MPORT_748_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_749_en & RAM_MPORT_749_mask) begin
      RAM[RAM_MPORT_749_addr] <= RAM_MPORT_749_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_750_en & RAM_MPORT_750_mask) begin
      RAM[RAM_MPORT_750_addr] <= RAM_MPORT_750_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_751_en & RAM_MPORT_751_mask) begin
      RAM[RAM_MPORT_751_addr] <= RAM_MPORT_751_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_752_en & RAM_MPORT_752_mask) begin
      RAM[RAM_MPORT_752_addr] <= RAM_MPORT_752_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_753_en & RAM_MPORT_753_mask) begin
      RAM[RAM_MPORT_753_addr] <= RAM_MPORT_753_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_754_en & RAM_MPORT_754_mask) begin
      RAM[RAM_MPORT_754_addr] <= RAM_MPORT_754_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_755_en & RAM_MPORT_755_mask) begin
      RAM[RAM_MPORT_755_addr] <= RAM_MPORT_755_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_756_en & RAM_MPORT_756_mask) begin
      RAM[RAM_MPORT_756_addr] <= RAM_MPORT_756_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_757_en & RAM_MPORT_757_mask) begin
      RAM[RAM_MPORT_757_addr] <= RAM_MPORT_757_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_758_en & RAM_MPORT_758_mask) begin
      RAM[RAM_MPORT_758_addr] <= RAM_MPORT_758_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_759_en & RAM_MPORT_759_mask) begin
      RAM[RAM_MPORT_759_addr] <= RAM_MPORT_759_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_760_en & RAM_MPORT_760_mask) begin
      RAM[RAM_MPORT_760_addr] <= RAM_MPORT_760_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_761_en & RAM_MPORT_761_mask) begin
      RAM[RAM_MPORT_761_addr] <= RAM_MPORT_761_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_762_en & RAM_MPORT_762_mask) begin
      RAM[RAM_MPORT_762_addr] <= RAM_MPORT_762_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_763_en & RAM_MPORT_763_mask) begin
      RAM[RAM_MPORT_763_addr] <= RAM_MPORT_763_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_764_en & RAM_MPORT_764_mask) begin
      RAM[RAM_MPORT_764_addr] <= RAM_MPORT_764_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_765_en & RAM_MPORT_765_mask) begin
      RAM[RAM_MPORT_765_addr] <= RAM_MPORT_765_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_766_en & RAM_MPORT_766_mask) begin
      RAM[RAM_MPORT_766_addr] <= RAM_MPORT_766_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_767_en & RAM_MPORT_767_mask) begin
      RAM[RAM_MPORT_767_addr] <= RAM_MPORT_767_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_768_en & RAM_MPORT_768_mask) begin
      RAM[RAM_MPORT_768_addr] <= RAM_MPORT_768_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_769_en & RAM_MPORT_769_mask) begin
      RAM[RAM_MPORT_769_addr] <= RAM_MPORT_769_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_770_en & RAM_MPORT_770_mask) begin
      RAM[RAM_MPORT_770_addr] <= RAM_MPORT_770_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_771_en & RAM_MPORT_771_mask) begin
      RAM[RAM_MPORT_771_addr] <= RAM_MPORT_771_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_772_en & RAM_MPORT_772_mask) begin
      RAM[RAM_MPORT_772_addr] <= RAM_MPORT_772_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_773_en & RAM_MPORT_773_mask) begin
      RAM[RAM_MPORT_773_addr] <= RAM_MPORT_773_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_774_en & RAM_MPORT_774_mask) begin
      RAM[RAM_MPORT_774_addr] <= RAM_MPORT_774_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_775_en & RAM_MPORT_775_mask) begin
      RAM[RAM_MPORT_775_addr] <= RAM_MPORT_775_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_776_en & RAM_MPORT_776_mask) begin
      RAM[RAM_MPORT_776_addr] <= RAM_MPORT_776_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_777_en & RAM_MPORT_777_mask) begin
      RAM[RAM_MPORT_777_addr] <= RAM_MPORT_777_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_778_en & RAM_MPORT_778_mask) begin
      RAM[RAM_MPORT_778_addr] <= RAM_MPORT_778_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_779_en & RAM_MPORT_779_mask) begin
      RAM[RAM_MPORT_779_addr] <= RAM_MPORT_779_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_780_en & RAM_MPORT_780_mask) begin
      RAM[RAM_MPORT_780_addr] <= RAM_MPORT_780_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_781_en & RAM_MPORT_781_mask) begin
      RAM[RAM_MPORT_781_addr] <= RAM_MPORT_781_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_782_en & RAM_MPORT_782_mask) begin
      RAM[RAM_MPORT_782_addr] <= RAM_MPORT_782_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_783_en & RAM_MPORT_783_mask) begin
      RAM[RAM_MPORT_783_addr] <= RAM_MPORT_783_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_784_en & RAM_MPORT_784_mask) begin
      RAM[RAM_MPORT_784_addr] <= RAM_MPORT_784_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_785_en & RAM_MPORT_785_mask) begin
      RAM[RAM_MPORT_785_addr] <= RAM_MPORT_785_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_786_en & RAM_MPORT_786_mask) begin
      RAM[RAM_MPORT_786_addr] <= RAM_MPORT_786_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_787_en & RAM_MPORT_787_mask) begin
      RAM[RAM_MPORT_787_addr] <= RAM_MPORT_787_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_788_en & RAM_MPORT_788_mask) begin
      RAM[RAM_MPORT_788_addr] <= RAM_MPORT_788_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_789_en & RAM_MPORT_789_mask) begin
      RAM[RAM_MPORT_789_addr] <= RAM_MPORT_789_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_790_en & RAM_MPORT_790_mask) begin
      RAM[RAM_MPORT_790_addr] <= RAM_MPORT_790_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_791_en & RAM_MPORT_791_mask) begin
      RAM[RAM_MPORT_791_addr] <= RAM_MPORT_791_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_792_en & RAM_MPORT_792_mask) begin
      RAM[RAM_MPORT_792_addr] <= RAM_MPORT_792_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_793_en & RAM_MPORT_793_mask) begin
      RAM[RAM_MPORT_793_addr] <= RAM_MPORT_793_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_794_en & RAM_MPORT_794_mask) begin
      RAM[RAM_MPORT_794_addr] <= RAM_MPORT_794_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_795_en & RAM_MPORT_795_mask) begin
      RAM[RAM_MPORT_795_addr] <= RAM_MPORT_795_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_796_en & RAM_MPORT_796_mask) begin
      RAM[RAM_MPORT_796_addr] <= RAM_MPORT_796_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_797_en & RAM_MPORT_797_mask) begin
      RAM[RAM_MPORT_797_addr] <= RAM_MPORT_797_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_798_en & RAM_MPORT_798_mask) begin
      RAM[RAM_MPORT_798_addr] <= RAM_MPORT_798_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_799_en & RAM_MPORT_799_mask) begin
      RAM[RAM_MPORT_799_addr] <= RAM_MPORT_799_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_800_en & RAM_MPORT_800_mask) begin
      RAM[RAM_MPORT_800_addr] <= RAM_MPORT_800_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_801_en & RAM_MPORT_801_mask) begin
      RAM[RAM_MPORT_801_addr] <= RAM_MPORT_801_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_802_en & RAM_MPORT_802_mask) begin
      RAM[RAM_MPORT_802_addr] <= RAM_MPORT_802_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_803_en & RAM_MPORT_803_mask) begin
      RAM[RAM_MPORT_803_addr] <= RAM_MPORT_803_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_804_en & RAM_MPORT_804_mask) begin
      RAM[RAM_MPORT_804_addr] <= RAM_MPORT_804_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_805_en & RAM_MPORT_805_mask) begin
      RAM[RAM_MPORT_805_addr] <= RAM_MPORT_805_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_806_en & RAM_MPORT_806_mask) begin
      RAM[RAM_MPORT_806_addr] <= RAM_MPORT_806_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_807_en & RAM_MPORT_807_mask) begin
      RAM[RAM_MPORT_807_addr] <= RAM_MPORT_807_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_808_en & RAM_MPORT_808_mask) begin
      RAM[RAM_MPORT_808_addr] <= RAM_MPORT_808_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_809_en & RAM_MPORT_809_mask) begin
      RAM[RAM_MPORT_809_addr] <= RAM_MPORT_809_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_810_en & RAM_MPORT_810_mask) begin
      RAM[RAM_MPORT_810_addr] <= RAM_MPORT_810_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_811_en & RAM_MPORT_811_mask) begin
      RAM[RAM_MPORT_811_addr] <= RAM_MPORT_811_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_812_en & RAM_MPORT_812_mask) begin
      RAM[RAM_MPORT_812_addr] <= RAM_MPORT_812_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_813_en & RAM_MPORT_813_mask) begin
      RAM[RAM_MPORT_813_addr] <= RAM_MPORT_813_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_814_en & RAM_MPORT_814_mask) begin
      RAM[RAM_MPORT_814_addr] <= RAM_MPORT_814_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_815_en & RAM_MPORT_815_mask) begin
      RAM[RAM_MPORT_815_addr] <= RAM_MPORT_815_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_816_en & RAM_MPORT_816_mask) begin
      RAM[RAM_MPORT_816_addr] <= RAM_MPORT_816_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_817_en & RAM_MPORT_817_mask) begin
      RAM[RAM_MPORT_817_addr] <= RAM_MPORT_817_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_818_en & RAM_MPORT_818_mask) begin
      RAM[RAM_MPORT_818_addr] <= RAM_MPORT_818_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_819_en & RAM_MPORT_819_mask) begin
      RAM[RAM_MPORT_819_addr] <= RAM_MPORT_819_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_820_en & RAM_MPORT_820_mask) begin
      RAM[RAM_MPORT_820_addr] <= RAM_MPORT_820_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_821_en & RAM_MPORT_821_mask) begin
      RAM[RAM_MPORT_821_addr] <= RAM_MPORT_821_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_822_en & RAM_MPORT_822_mask) begin
      RAM[RAM_MPORT_822_addr] <= RAM_MPORT_822_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_823_en & RAM_MPORT_823_mask) begin
      RAM[RAM_MPORT_823_addr] <= RAM_MPORT_823_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_824_en & RAM_MPORT_824_mask) begin
      RAM[RAM_MPORT_824_addr] <= RAM_MPORT_824_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_825_en & RAM_MPORT_825_mask) begin
      RAM[RAM_MPORT_825_addr] <= RAM_MPORT_825_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_826_en & RAM_MPORT_826_mask) begin
      RAM[RAM_MPORT_826_addr] <= RAM_MPORT_826_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_827_en & RAM_MPORT_827_mask) begin
      RAM[RAM_MPORT_827_addr] <= RAM_MPORT_827_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_828_en & RAM_MPORT_828_mask) begin
      RAM[RAM_MPORT_828_addr] <= RAM_MPORT_828_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_829_en & RAM_MPORT_829_mask) begin
      RAM[RAM_MPORT_829_addr] <= RAM_MPORT_829_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_830_en & RAM_MPORT_830_mask) begin
      RAM[RAM_MPORT_830_addr] <= RAM_MPORT_830_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_831_en & RAM_MPORT_831_mask) begin
      RAM[RAM_MPORT_831_addr] <= RAM_MPORT_831_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_832_en & RAM_MPORT_832_mask) begin
      RAM[RAM_MPORT_832_addr] <= RAM_MPORT_832_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_833_en & RAM_MPORT_833_mask) begin
      RAM[RAM_MPORT_833_addr] <= RAM_MPORT_833_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_834_en & RAM_MPORT_834_mask) begin
      RAM[RAM_MPORT_834_addr] <= RAM_MPORT_834_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_835_en & RAM_MPORT_835_mask) begin
      RAM[RAM_MPORT_835_addr] <= RAM_MPORT_835_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_836_en & RAM_MPORT_836_mask) begin
      RAM[RAM_MPORT_836_addr] <= RAM_MPORT_836_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_837_en & RAM_MPORT_837_mask) begin
      RAM[RAM_MPORT_837_addr] <= RAM_MPORT_837_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_838_en & RAM_MPORT_838_mask) begin
      RAM[RAM_MPORT_838_addr] <= RAM_MPORT_838_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_839_en & RAM_MPORT_839_mask) begin
      RAM[RAM_MPORT_839_addr] <= RAM_MPORT_839_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_840_en & RAM_MPORT_840_mask) begin
      RAM[RAM_MPORT_840_addr] <= RAM_MPORT_840_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_841_en & RAM_MPORT_841_mask) begin
      RAM[RAM_MPORT_841_addr] <= RAM_MPORT_841_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_842_en & RAM_MPORT_842_mask) begin
      RAM[RAM_MPORT_842_addr] <= RAM_MPORT_842_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_843_en & RAM_MPORT_843_mask) begin
      RAM[RAM_MPORT_843_addr] <= RAM_MPORT_843_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_844_en & RAM_MPORT_844_mask) begin
      RAM[RAM_MPORT_844_addr] <= RAM_MPORT_844_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_845_en & RAM_MPORT_845_mask) begin
      RAM[RAM_MPORT_845_addr] <= RAM_MPORT_845_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_846_en & RAM_MPORT_846_mask) begin
      RAM[RAM_MPORT_846_addr] <= RAM_MPORT_846_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_847_en & RAM_MPORT_847_mask) begin
      RAM[RAM_MPORT_847_addr] <= RAM_MPORT_847_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_848_en & RAM_MPORT_848_mask) begin
      RAM[RAM_MPORT_848_addr] <= RAM_MPORT_848_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_849_en & RAM_MPORT_849_mask) begin
      RAM[RAM_MPORT_849_addr] <= RAM_MPORT_849_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_850_en & RAM_MPORT_850_mask) begin
      RAM[RAM_MPORT_850_addr] <= RAM_MPORT_850_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_851_en & RAM_MPORT_851_mask) begin
      RAM[RAM_MPORT_851_addr] <= RAM_MPORT_851_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_852_en & RAM_MPORT_852_mask) begin
      RAM[RAM_MPORT_852_addr] <= RAM_MPORT_852_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_853_en & RAM_MPORT_853_mask) begin
      RAM[RAM_MPORT_853_addr] <= RAM_MPORT_853_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_854_en & RAM_MPORT_854_mask) begin
      RAM[RAM_MPORT_854_addr] <= RAM_MPORT_854_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_855_en & RAM_MPORT_855_mask) begin
      RAM[RAM_MPORT_855_addr] <= RAM_MPORT_855_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_856_en & RAM_MPORT_856_mask) begin
      RAM[RAM_MPORT_856_addr] <= RAM_MPORT_856_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_857_en & RAM_MPORT_857_mask) begin
      RAM[RAM_MPORT_857_addr] <= RAM_MPORT_857_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_858_en & RAM_MPORT_858_mask) begin
      RAM[RAM_MPORT_858_addr] <= RAM_MPORT_858_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_859_en & RAM_MPORT_859_mask) begin
      RAM[RAM_MPORT_859_addr] <= RAM_MPORT_859_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_860_en & RAM_MPORT_860_mask) begin
      RAM[RAM_MPORT_860_addr] <= RAM_MPORT_860_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_861_en & RAM_MPORT_861_mask) begin
      RAM[RAM_MPORT_861_addr] <= RAM_MPORT_861_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_862_en & RAM_MPORT_862_mask) begin
      RAM[RAM_MPORT_862_addr] <= RAM_MPORT_862_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_863_en & RAM_MPORT_863_mask) begin
      RAM[RAM_MPORT_863_addr] <= RAM_MPORT_863_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_864_en & RAM_MPORT_864_mask) begin
      RAM[RAM_MPORT_864_addr] <= RAM_MPORT_864_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_865_en & RAM_MPORT_865_mask) begin
      RAM[RAM_MPORT_865_addr] <= RAM_MPORT_865_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_866_en & RAM_MPORT_866_mask) begin
      RAM[RAM_MPORT_866_addr] <= RAM_MPORT_866_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_867_en & RAM_MPORT_867_mask) begin
      RAM[RAM_MPORT_867_addr] <= RAM_MPORT_867_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_868_en & RAM_MPORT_868_mask) begin
      RAM[RAM_MPORT_868_addr] <= RAM_MPORT_868_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_869_en & RAM_MPORT_869_mask) begin
      RAM[RAM_MPORT_869_addr] <= RAM_MPORT_869_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_870_en & RAM_MPORT_870_mask) begin
      RAM[RAM_MPORT_870_addr] <= RAM_MPORT_870_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_871_en & RAM_MPORT_871_mask) begin
      RAM[RAM_MPORT_871_addr] <= RAM_MPORT_871_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_872_en & RAM_MPORT_872_mask) begin
      RAM[RAM_MPORT_872_addr] <= RAM_MPORT_872_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_873_en & RAM_MPORT_873_mask) begin
      RAM[RAM_MPORT_873_addr] <= RAM_MPORT_873_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_874_en & RAM_MPORT_874_mask) begin
      RAM[RAM_MPORT_874_addr] <= RAM_MPORT_874_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_875_en & RAM_MPORT_875_mask) begin
      RAM[RAM_MPORT_875_addr] <= RAM_MPORT_875_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_876_en & RAM_MPORT_876_mask) begin
      RAM[RAM_MPORT_876_addr] <= RAM_MPORT_876_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_877_en & RAM_MPORT_877_mask) begin
      RAM[RAM_MPORT_877_addr] <= RAM_MPORT_877_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_878_en & RAM_MPORT_878_mask) begin
      RAM[RAM_MPORT_878_addr] <= RAM_MPORT_878_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_879_en & RAM_MPORT_879_mask) begin
      RAM[RAM_MPORT_879_addr] <= RAM_MPORT_879_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_880_en & RAM_MPORT_880_mask) begin
      RAM[RAM_MPORT_880_addr] <= RAM_MPORT_880_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_881_en & RAM_MPORT_881_mask) begin
      RAM[RAM_MPORT_881_addr] <= RAM_MPORT_881_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_882_en & RAM_MPORT_882_mask) begin
      RAM[RAM_MPORT_882_addr] <= RAM_MPORT_882_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_883_en & RAM_MPORT_883_mask) begin
      RAM[RAM_MPORT_883_addr] <= RAM_MPORT_883_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_884_en & RAM_MPORT_884_mask) begin
      RAM[RAM_MPORT_884_addr] <= RAM_MPORT_884_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_885_en & RAM_MPORT_885_mask) begin
      RAM[RAM_MPORT_885_addr] <= RAM_MPORT_885_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_886_en & RAM_MPORT_886_mask) begin
      RAM[RAM_MPORT_886_addr] <= RAM_MPORT_886_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_887_en & RAM_MPORT_887_mask) begin
      RAM[RAM_MPORT_887_addr] <= RAM_MPORT_887_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_888_en & RAM_MPORT_888_mask) begin
      RAM[RAM_MPORT_888_addr] <= RAM_MPORT_888_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_889_en & RAM_MPORT_889_mask) begin
      RAM[RAM_MPORT_889_addr] <= RAM_MPORT_889_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_890_en & RAM_MPORT_890_mask) begin
      RAM[RAM_MPORT_890_addr] <= RAM_MPORT_890_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_891_en & RAM_MPORT_891_mask) begin
      RAM[RAM_MPORT_891_addr] <= RAM_MPORT_891_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_892_en & RAM_MPORT_892_mask) begin
      RAM[RAM_MPORT_892_addr] <= RAM_MPORT_892_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_893_en & RAM_MPORT_893_mask) begin
      RAM[RAM_MPORT_893_addr] <= RAM_MPORT_893_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_894_en & RAM_MPORT_894_mask) begin
      RAM[RAM_MPORT_894_addr] <= RAM_MPORT_894_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_895_en & RAM_MPORT_895_mask) begin
      RAM[RAM_MPORT_895_addr] <= RAM_MPORT_895_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_896_en & RAM_MPORT_896_mask) begin
      RAM[RAM_MPORT_896_addr] <= RAM_MPORT_896_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_897_en & RAM_MPORT_897_mask) begin
      RAM[RAM_MPORT_897_addr] <= RAM_MPORT_897_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_898_en & RAM_MPORT_898_mask) begin
      RAM[RAM_MPORT_898_addr] <= RAM_MPORT_898_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_899_en & RAM_MPORT_899_mask) begin
      RAM[RAM_MPORT_899_addr] <= RAM_MPORT_899_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_900_en & RAM_MPORT_900_mask) begin
      RAM[RAM_MPORT_900_addr] <= RAM_MPORT_900_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_901_en & RAM_MPORT_901_mask) begin
      RAM[RAM_MPORT_901_addr] <= RAM_MPORT_901_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_902_en & RAM_MPORT_902_mask) begin
      RAM[RAM_MPORT_902_addr] <= RAM_MPORT_902_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_903_en & RAM_MPORT_903_mask) begin
      RAM[RAM_MPORT_903_addr] <= RAM_MPORT_903_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_904_en & RAM_MPORT_904_mask) begin
      RAM[RAM_MPORT_904_addr] <= RAM_MPORT_904_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_905_en & RAM_MPORT_905_mask) begin
      RAM[RAM_MPORT_905_addr] <= RAM_MPORT_905_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_906_en & RAM_MPORT_906_mask) begin
      RAM[RAM_MPORT_906_addr] <= RAM_MPORT_906_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_907_en & RAM_MPORT_907_mask) begin
      RAM[RAM_MPORT_907_addr] <= RAM_MPORT_907_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_908_en & RAM_MPORT_908_mask) begin
      RAM[RAM_MPORT_908_addr] <= RAM_MPORT_908_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_909_en & RAM_MPORT_909_mask) begin
      RAM[RAM_MPORT_909_addr] <= RAM_MPORT_909_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_910_en & RAM_MPORT_910_mask) begin
      RAM[RAM_MPORT_910_addr] <= RAM_MPORT_910_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_911_en & RAM_MPORT_911_mask) begin
      RAM[RAM_MPORT_911_addr] <= RAM_MPORT_911_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_912_en & RAM_MPORT_912_mask) begin
      RAM[RAM_MPORT_912_addr] <= RAM_MPORT_912_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_913_en & RAM_MPORT_913_mask) begin
      RAM[RAM_MPORT_913_addr] <= RAM_MPORT_913_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_914_en & RAM_MPORT_914_mask) begin
      RAM[RAM_MPORT_914_addr] <= RAM_MPORT_914_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_915_en & RAM_MPORT_915_mask) begin
      RAM[RAM_MPORT_915_addr] <= RAM_MPORT_915_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_916_en & RAM_MPORT_916_mask) begin
      RAM[RAM_MPORT_916_addr] <= RAM_MPORT_916_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_917_en & RAM_MPORT_917_mask) begin
      RAM[RAM_MPORT_917_addr] <= RAM_MPORT_917_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_918_en & RAM_MPORT_918_mask) begin
      RAM[RAM_MPORT_918_addr] <= RAM_MPORT_918_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_919_en & RAM_MPORT_919_mask) begin
      RAM[RAM_MPORT_919_addr] <= RAM_MPORT_919_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_920_en & RAM_MPORT_920_mask) begin
      RAM[RAM_MPORT_920_addr] <= RAM_MPORT_920_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_921_en & RAM_MPORT_921_mask) begin
      RAM[RAM_MPORT_921_addr] <= RAM_MPORT_921_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_922_en & RAM_MPORT_922_mask) begin
      RAM[RAM_MPORT_922_addr] <= RAM_MPORT_922_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_923_en & RAM_MPORT_923_mask) begin
      RAM[RAM_MPORT_923_addr] <= RAM_MPORT_923_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_924_en & RAM_MPORT_924_mask) begin
      RAM[RAM_MPORT_924_addr] <= RAM_MPORT_924_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_925_en & RAM_MPORT_925_mask) begin
      RAM[RAM_MPORT_925_addr] <= RAM_MPORT_925_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_926_en & RAM_MPORT_926_mask) begin
      RAM[RAM_MPORT_926_addr] <= RAM_MPORT_926_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_927_en & RAM_MPORT_927_mask) begin
      RAM[RAM_MPORT_927_addr] <= RAM_MPORT_927_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_928_en & RAM_MPORT_928_mask) begin
      RAM[RAM_MPORT_928_addr] <= RAM_MPORT_928_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_929_en & RAM_MPORT_929_mask) begin
      RAM[RAM_MPORT_929_addr] <= RAM_MPORT_929_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_930_en & RAM_MPORT_930_mask) begin
      RAM[RAM_MPORT_930_addr] <= RAM_MPORT_930_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_931_en & RAM_MPORT_931_mask) begin
      RAM[RAM_MPORT_931_addr] <= RAM_MPORT_931_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_932_en & RAM_MPORT_932_mask) begin
      RAM[RAM_MPORT_932_addr] <= RAM_MPORT_932_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_933_en & RAM_MPORT_933_mask) begin
      RAM[RAM_MPORT_933_addr] <= RAM_MPORT_933_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_934_en & RAM_MPORT_934_mask) begin
      RAM[RAM_MPORT_934_addr] <= RAM_MPORT_934_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_935_en & RAM_MPORT_935_mask) begin
      RAM[RAM_MPORT_935_addr] <= RAM_MPORT_935_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_936_en & RAM_MPORT_936_mask) begin
      RAM[RAM_MPORT_936_addr] <= RAM_MPORT_936_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_937_en & RAM_MPORT_937_mask) begin
      RAM[RAM_MPORT_937_addr] <= RAM_MPORT_937_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_938_en & RAM_MPORT_938_mask) begin
      RAM[RAM_MPORT_938_addr] <= RAM_MPORT_938_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_939_en & RAM_MPORT_939_mask) begin
      RAM[RAM_MPORT_939_addr] <= RAM_MPORT_939_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_940_en & RAM_MPORT_940_mask) begin
      RAM[RAM_MPORT_940_addr] <= RAM_MPORT_940_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_941_en & RAM_MPORT_941_mask) begin
      RAM[RAM_MPORT_941_addr] <= RAM_MPORT_941_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_942_en & RAM_MPORT_942_mask) begin
      RAM[RAM_MPORT_942_addr] <= RAM_MPORT_942_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_943_en & RAM_MPORT_943_mask) begin
      RAM[RAM_MPORT_943_addr] <= RAM_MPORT_943_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_944_en & RAM_MPORT_944_mask) begin
      RAM[RAM_MPORT_944_addr] <= RAM_MPORT_944_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_945_en & RAM_MPORT_945_mask) begin
      RAM[RAM_MPORT_945_addr] <= RAM_MPORT_945_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_946_en & RAM_MPORT_946_mask) begin
      RAM[RAM_MPORT_946_addr] <= RAM_MPORT_946_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_947_en & RAM_MPORT_947_mask) begin
      RAM[RAM_MPORT_947_addr] <= RAM_MPORT_947_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_948_en & RAM_MPORT_948_mask) begin
      RAM[RAM_MPORT_948_addr] <= RAM_MPORT_948_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_949_en & RAM_MPORT_949_mask) begin
      RAM[RAM_MPORT_949_addr] <= RAM_MPORT_949_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_950_en & RAM_MPORT_950_mask) begin
      RAM[RAM_MPORT_950_addr] <= RAM_MPORT_950_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_951_en & RAM_MPORT_951_mask) begin
      RAM[RAM_MPORT_951_addr] <= RAM_MPORT_951_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_952_en & RAM_MPORT_952_mask) begin
      RAM[RAM_MPORT_952_addr] <= RAM_MPORT_952_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_953_en & RAM_MPORT_953_mask) begin
      RAM[RAM_MPORT_953_addr] <= RAM_MPORT_953_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_954_en & RAM_MPORT_954_mask) begin
      RAM[RAM_MPORT_954_addr] <= RAM_MPORT_954_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_955_en & RAM_MPORT_955_mask) begin
      RAM[RAM_MPORT_955_addr] <= RAM_MPORT_955_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_956_en & RAM_MPORT_956_mask) begin
      RAM[RAM_MPORT_956_addr] <= RAM_MPORT_956_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_957_en & RAM_MPORT_957_mask) begin
      RAM[RAM_MPORT_957_addr] <= RAM_MPORT_957_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_958_en & RAM_MPORT_958_mask) begin
      RAM[RAM_MPORT_958_addr] <= RAM_MPORT_958_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_959_en & RAM_MPORT_959_mask) begin
      RAM[RAM_MPORT_959_addr] <= RAM_MPORT_959_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_960_en & RAM_MPORT_960_mask) begin
      RAM[RAM_MPORT_960_addr] <= RAM_MPORT_960_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_961_en & RAM_MPORT_961_mask) begin
      RAM[RAM_MPORT_961_addr] <= RAM_MPORT_961_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_962_en & RAM_MPORT_962_mask) begin
      RAM[RAM_MPORT_962_addr] <= RAM_MPORT_962_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_963_en & RAM_MPORT_963_mask) begin
      RAM[RAM_MPORT_963_addr] <= RAM_MPORT_963_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_964_en & RAM_MPORT_964_mask) begin
      RAM[RAM_MPORT_964_addr] <= RAM_MPORT_964_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_965_en & RAM_MPORT_965_mask) begin
      RAM[RAM_MPORT_965_addr] <= RAM_MPORT_965_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_966_en & RAM_MPORT_966_mask) begin
      RAM[RAM_MPORT_966_addr] <= RAM_MPORT_966_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_967_en & RAM_MPORT_967_mask) begin
      RAM[RAM_MPORT_967_addr] <= RAM_MPORT_967_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_968_en & RAM_MPORT_968_mask) begin
      RAM[RAM_MPORT_968_addr] <= RAM_MPORT_968_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_969_en & RAM_MPORT_969_mask) begin
      RAM[RAM_MPORT_969_addr] <= RAM_MPORT_969_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_970_en & RAM_MPORT_970_mask) begin
      RAM[RAM_MPORT_970_addr] <= RAM_MPORT_970_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_971_en & RAM_MPORT_971_mask) begin
      RAM[RAM_MPORT_971_addr] <= RAM_MPORT_971_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_972_en & RAM_MPORT_972_mask) begin
      RAM[RAM_MPORT_972_addr] <= RAM_MPORT_972_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_973_en & RAM_MPORT_973_mask) begin
      RAM[RAM_MPORT_973_addr] <= RAM_MPORT_973_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_974_en & RAM_MPORT_974_mask) begin
      RAM[RAM_MPORT_974_addr] <= RAM_MPORT_974_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_975_en & RAM_MPORT_975_mask) begin
      RAM[RAM_MPORT_975_addr] <= RAM_MPORT_975_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_976_en & RAM_MPORT_976_mask) begin
      RAM[RAM_MPORT_976_addr] <= RAM_MPORT_976_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_977_en & RAM_MPORT_977_mask) begin
      RAM[RAM_MPORT_977_addr] <= RAM_MPORT_977_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_978_en & RAM_MPORT_978_mask) begin
      RAM[RAM_MPORT_978_addr] <= RAM_MPORT_978_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_979_en & RAM_MPORT_979_mask) begin
      RAM[RAM_MPORT_979_addr] <= RAM_MPORT_979_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_980_en & RAM_MPORT_980_mask) begin
      RAM[RAM_MPORT_980_addr] <= RAM_MPORT_980_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_981_en & RAM_MPORT_981_mask) begin
      RAM[RAM_MPORT_981_addr] <= RAM_MPORT_981_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_982_en & RAM_MPORT_982_mask) begin
      RAM[RAM_MPORT_982_addr] <= RAM_MPORT_982_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_983_en & RAM_MPORT_983_mask) begin
      RAM[RAM_MPORT_983_addr] <= RAM_MPORT_983_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_984_en & RAM_MPORT_984_mask) begin
      RAM[RAM_MPORT_984_addr] <= RAM_MPORT_984_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_985_en & RAM_MPORT_985_mask) begin
      RAM[RAM_MPORT_985_addr] <= RAM_MPORT_985_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_986_en & RAM_MPORT_986_mask) begin
      RAM[RAM_MPORT_986_addr] <= RAM_MPORT_986_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_987_en & RAM_MPORT_987_mask) begin
      RAM[RAM_MPORT_987_addr] <= RAM_MPORT_987_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_988_en & RAM_MPORT_988_mask) begin
      RAM[RAM_MPORT_988_addr] <= RAM_MPORT_988_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_989_en & RAM_MPORT_989_mask) begin
      RAM[RAM_MPORT_989_addr] <= RAM_MPORT_989_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_990_en & RAM_MPORT_990_mask) begin
      RAM[RAM_MPORT_990_addr] <= RAM_MPORT_990_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_991_en & RAM_MPORT_991_mask) begin
      RAM[RAM_MPORT_991_addr] <= RAM_MPORT_991_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_992_en & RAM_MPORT_992_mask) begin
      RAM[RAM_MPORT_992_addr] <= RAM_MPORT_992_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_993_en & RAM_MPORT_993_mask) begin
      RAM[RAM_MPORT_993_addr] <= RAM_MPORT_993_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_994_en & RAM_MPORT_994_mask) begin
      RAM[RAM_MPORT_994_addr] <= RAM_MPORT_994_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_995_en & RAM_MPORT_995_mask) begin
      RAM[RAM_MPORT_995_addr] <= RAM_MPORT_995_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_996_en & RAM_MPORT_996_mask) begin
      RAM[RAM_MPORT_996_addr] <= RAM_MPORT_996_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_997_en & RAM_MPORT_997_mask) begin
      RAM[RAM_MPORT_997_addr] <= RAM_MPORT_997_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_998_en & RAM_MPORT_998_mask) begin
      RAM[RAM_MPORT_998_addr] <= RAM_MPORT_998_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_999_en & RAM_MPORT_999_mask) begin
      RAM[RAM_MPORT_999_addr] <= RAM_MPORT_999_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1000_en & RAM_MPORT_1000_mask) begin
      RAM[RAM_MPORT_1000_addr] <= RAM_MPORT_1000_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1001_en & RAM_MPORT_1001_mask) begin
      RAM[RAM_MPORT_1001_addr] <= RAM_MPORT_1001_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1002_en & RAM_MPORT_1002_mask) begin
      RAM[RAM_MPORT_1002_addr] <= RAM_MPORT_1002_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1003_en & RAM_MPORT_1003_mask) begin
      RAM[RAM_MPORT_1003_addr] <= RAM_MPORT_1003_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1004_en & RAM_MPORT_1004_mask) begin
      RAM[RAM_MPORT_1004_addr] <= RAM_MPORT_1004_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1005_en & RAM_MPORT_1005_mask) begin
      RAM[RAM_MPORT_1005_addr] <= RAM_MPORT_1005_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1006_en & RAM_MPORT_1006_mask) begin
      RAM[RAM_MPORT_1006_addr] <= RAM_MPORT_1006_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1007_en & RAM_MPORT_1007_mask) begin
      RAM[RAM_MPORT_1007_addr] <= RAM_MPORT_1007_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1008_en & RAM_MPORT_1008_mask) begin
      RAM[RAM_MPORT_1008_addr] <= RAM_MPORT_1008_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1009_en & RAM_MPORT_1009_mask) begin
      RAM[RAM_MPORT_1009_addr] <= RAM_MPORT_1009_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1010_en & RAM_MPORT_1010_mask) begin
      RAM[RAM_MPORT_1010_addr] <= RAM_MPORT_1010_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1011_en & RAM_MPORT_1011_mask) begin
      RAM[RAM_MPORT_1011_addr] <= RAM_MPORT_1011_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1012_en & RAM_MPORT_1012_mask) begin
      RAM[RAM_MPORT_1012_addr] <= RAM_MPORT_1012_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1013_en & RAM_MPORT_1013_mask) begin
      RAM[RAM_MPORT_1013_addr] <= RAM_MPORT_1013_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1014_en & RAM_MPORT_1014_mask) begin
      RAM[RAM_MPORT_1014_addr] <= RAM_MPORT_1014_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1015_en & RAM_MPORT_1015_mask) begin
      RAM[RAM_MPORT_1015_addr] <= RAM_MPORT_1015_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1016_en & RAM_MPORT_1016_mask) begin
      RAM[RAM_MPORT_1016_addr] <= RAM_MPORT_1016_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1017_en & RAM_MPORT_1017_mask) begin
      RAM[RAM_MPORT_1017_addr] <= RAM_MPORT_1017_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1018_en & RAM_MPORT_1018_mask) begin
      RAM[RAM_MPORT_1018_addr] <= RAM_MPORT_1018_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1019_en & RAM_MPORT_1019_mask) begin
      RAM[RAM_MPORT_1019_addr] <= RAM_MPORT_1019_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1020_en & RAM_MPORT_1020_mask) begin
      RAM[RAM_MPORT_1020_addr] <= RAM_MPORT_1020_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1021_en & RAM_MPORT_1021_mask) begin
      RAM[RAM_MPORT_1021_addr] <= RAM_MPORT_1021_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1022_en & RAM_MPORT_1022_mask) begin
      RAM[RAM_MPORT_1022_addr] <= RAM_MPORT_1022_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1023_en & RAM_MPORT_1023_mask) begin
      RAM[RAM_MPORT_1023_addr] <= RAM_MPORT_1023_data; // @[DM.scala 12:29]
    end
    if (RAM_MPORT_1024_en & RAM_MPORT_1024_mask) begin
      RAM[RAM_MPORT_1024_addr] <= RAM_MPORT_1024_data; // @[DM.scala 12:29]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & io_WE & ~reset) begin
          $fwrite(32'h80000002,"@0x%x: 0x%x <= 0x%x\n",io_PC,io_Addr,io_WD); // @[DM.scala 21:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    RAM[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EXT(
  input  [15:0] io_imm16,
  input         io_IsSignEXT,
  output [31:0] io_imm32
);
  wire [31:0] _io_imm32_T = {16'hffff,io_imm16}; // @[Cat.scala 31:58]
  wire [31:0] _io_imm32_T_1 = {16'h0,io_imm16}; // @[Cat.scala 31:58]
  assign io_imm32 = io_IsSignEXT & io_imm16[15] ? _io_imm32_T : _io_imm32_T_1; // @[EXT.scala 12:57 13:18 15:18]
endmodule
module DataPath(
  input         clock,
  input         reset,
  input         io_WEGRF,
  input         io_WEDM,
  input  [1:0]  io_RegDst,
  input  [1:0]  io_WhichToReg,
  input  [3:0]  io_ALUOp,
  input         io_ALUSrc,
  input         io_IsSignExt,
  input         io_IsBranchType,
  input         io_IsJType,
  input         io_IsJr,
  output [31:0] io_instr,
  output        io_IsEq
);
  wire  IFU_Module_clock; // @[DataPath.scala 21:33]
  wire  IFU_Module_reset; // @[DataPath.scala 21:33]
  wire [31:0] IFU_Module_io_NPC; // @[DataPath.scala 21:33]
  wire [31:0] IFU_Module_io_instr; // @[DataPath.scala 21:33]
  wire [31:0] IFU_Module_io_PC; // @[DataPath.scala 21:33]
  wire [31:0] NPC_Module_io_PC; // @[DataPath.scala 22:33]
  wire  NPC_Module_io_IsBranchType; // @[DataPath.scala 22:33]
  wire  NPC_Module_io_IsJType; // @[DataPath.scala 22:33]
  wire [31:0] NPC_Module_io_instr; // @[DataPath.scala 22:33]
  wire  NPC_Module_io_IsJr; // @[DataPath.scala 22:33]
  wire [31:0] NPC_Module_io_JrAddr; // @[DataPath.scala 22:33]
  wire [31:0] NPC_Module_io_imm32; // @[DataPath.scala 22:33]
  wire [31:0] NPC_Module_io_NPC; // @[DataPath.scala 22:33]
  wire  GRF_Module_clock; // @[DataPath.scala 23:33]
  wire  GRF_Module_reset; // @[DataPath.scala 23:33]
  wire [4:0] GRF_Module_io_A1; // @[DataPath.scala 23:33]
  wire [4:0] GRF_Module_io_A2; // @[DataPath.scala 23:33]
  wire [4:0] GRF_Module_io_A3; // @[DataPath.scala 23:33]
  wire  GRF_Module_io_WE; // @[DataPath.scala 23:33]
  wire [31:0] GRF_Module_io_WD; // @[DataPath.scala 23:33]
  wire [31:0] GRF_Module_io_PC; // @[DataPath.scala 23:33]
  wire [31:0] GRF_Module_io_O1; // @[DataPath.scala 23:33]
  wire [31:0] GRF_Module_io_O2; // @[DataPath.scala 23:33]
  wire [31:0] ALU_Module_io_A1; // @[DataPath.scala 24:33]
  wire [31:0] ALU_Module_io_A2; // @[DataPath.scala 24:33]
  wire [3:0] ALU_Module_io_ALUOp; // @[DataPath.scala 24:33]
  wire [31:0] ALU_Module_io_O; // @[DataPath.scala 24:33]
  wire  ALU_Module_io_IsEq; // @[DataPath.scala 24:33]
  wire  DM_Module_clock; // @[DataPath.scala 25:31]
  wire  DM_Module_reset; // @[DataPath.scala 25:31]
  wire [31:0] DM_Module_io_Addr; // @[DataPath.scala 25:31]
  wire [31:0] DM_Module_io_WD; // @[DataPath.scala 25:31]
  wire  DM_Module_io_WE; // @[DataPath.scala 25:31]
  wire [31:0] DM_Module_io_PC; // @[DataPath.scala 25:31]
  wire [31:0] DM_Module_io_RD; // @[DataPath.scala 25:31]
  wire [15:0] EXT_Module_io_imm16; // @[DataPath.scala 26:33]
  wire  EXT_Module_io_IsSignEXT; // @[DataPath.scala 26:33]
  wire [31:0] EXT_Module_io_imm32; // @[DataPath.scala 26:33]
  wire  _GRFWriteAddr_T = io_RegDst == 2'h0; // @[DataPath.scala 38:60]
  wire  _GRFWriteAddr_T_2 = io_RegDst == 2'h1; // @[DataPath.scala 39:59]
  wire  _GRFWriteAddr_T_4 = io_RegDst == 2'h2; // @[DataPath.scala 40:59]
  wire [4:0] _GRFWriteAddr_T_5 = _GRFWriteAddr_T_4 ? 5'h1f : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _GRFWriteAddr_T_6 = _GRFWriteAddr_T_2 ? IFU_Module_io_instr[20:16] : _GRFWriteAddr_T_5; // @[Mux.scala 101:16]
  wire  _GRFWrite_T = io_WhichToReg == 2'h0; // @[DataPath.scala 41:60]
  wire  _GRFWrite_T_1 = io_WhichToReg == 2'h1; // @[DataPath.scala 42:60]
  wire  _GRFWrite_T_2 = io_WhichToReg == 2'h2; // @[DataPath.scala 43:60]
  wire [31:0] _GRFWrite_T_4 = IFU_Module_io_PC + 32'h4; // @[DataPath.scala 43:90]
  wire [31:0] _GRFWrite_T_5 = _GRFWrite_T_2 ? _GRFWrite_T_4 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _GRFWrite_T_6 = _GRFWrite_T_1 ? DM_Module_io_RD : _GRFWrite_T_5; // @[Mux.scala 101:16]
  wire  _ALURead2_T = ~io_ALUSrc; // @[DataPath.scala 52:56]
  wire [31:0] _ALURead2_T_2 = io_ALUSrc ? EXT_Module_io_imm32 : 32'h0; // @[Mux.scala 101:16]
  IFU IFU_Module ( // @[DataPath.scala 21:33]
    .clock(IFU_Module_clock),
    .reset(IFU_Module_reset),
    .io_NPC(IFU_Module_io_NPC),
    .io_instr(IFU_Module_io_instr),
    .io_PC(IFU_Module_io_PC)
  );
  NPC NPC_Module ( // @[DataPath.scala 22:33]
    .io_PC(NPC_Module_io_PC),
    .io_IsBranchType(NPC_Module_io_IsBranchType),
    .io_IsJType(NPC_Module_io_IsJType),
    .io_instr(NPC_Module_io_instr),
    .io_IsJr(NPC_Module_io_IsJr),
    .io_JrAddr(NPC_Module_io_JrAddr),
    .io_imm32(NPC_Module_io_imm32),
    .io_NPC(NPC_Module_io_NPC)
  );
  GRF GRF_Module ( // @[DataPath.scala 23:33]
    .clock(GRF_Module_clock),
    .reset(GRF_Module_reset),
    .io_A1(GRF_Module_io_A1),
    .io_A2(GRF_Module_io_A2),
    .io_A3(GRF_Module_io_A3),
    .io_WE(GRF_Module_io_WE),
    .io_WD(GRF_Module_io_WD),
    .io_PC(GRF_Module_io_PC),
    .io_O1(GRF_Module_io_O1),
    .io_O2(GRF_Module_io_O2)
  );
  ALU ALU_Module ( // @[DataPath.scala 24:33]
    .io_A1(ALU_Module_io_A1),
    .io_A2(ALU_Module_io_A2),
    .io_ALUOp(ALU_Module_io_ALUOp),
    .io_O(ALU_Module_io_O),
    .io_IsEq(ALU_Module_io_IsEq)
  );
  DM DM_Module ( // @[DataPath.scala 25:31]
    .clock(DM_Module_clock),
    .reset(DM_Module_reset),
    .io_Addr(DM_Module_io_Addr),
    .io_WD(DM_Module_io_WD),
    .io_WE(DM_Module_io_WE),
    .io_PC(DM_Module_io_PC),
    .io_RD(DM_Module_io_RD)
  );
  EXT EXT_Module ( // @[DataPath.scala 26:33]
    .io_imm16(EXT_Module_io_imm16),
    .io_IsSignEXT(EXT_Module_io_IsSignEXT),
    .io_imm32(EXT_Module_io_imm32)
  );
  assign io_instr = IFU_Module_io_instr; // @[DataPath.scala 67:14]
  assign io_IsEq = ALU_Module_io_IsEq; // @[DataPath.scala 68:13]
  assign IFU_Module_clock = clock;
  assign IFU_Module_reset = reset;
  assign IFU_Module_io_NPC = NPC_Module_io_NPC; // @[DataPath.scala 28:23]
  assign NPC_Module_io_PC = IFU_Module_io_PC; // @[DataPath.scala 30:22]
  assign NPC_Module_io_IsBranchType = io_IsBranchType; // @[DataPath.scala 31:32]
  assign NPC_Module_io_IsJType = io_IsJType; // @[DataPath.scala 32:27]
  assign NPC_Module_io_instr = IFU_Module_io_instr; // @[DataPath.scala 33:25]
  assign NPC_Module_io_IsJr = io_IsJr; // @[DataPath.scala 34:24]
  assign NPC_Module_io_JrAddr = GRF_Module_io_O1; // @[DataPath.scala 35:26]
  assign NPC_Module_io_imm32 = EXT_Module_io_imm32; // @[DataPath.scala 36:25]
  assign GRF_Module_clock = clock;
  assign GRF_Module_reset = reset;
  assign GRF_Module_io_A1 = IFU_Module_io_instr[25:21]; // @[DataPath.scala 45:44]
  assign GRF_Module_io_A2 = IFU_Module_io_instr[20:16]; // @[DataPath.scala 46:44]
  assign GRF_Module_io_A3 = _GRFWriteAddr_T ? IFU_Module_io_instr[15:11] : _GRFWriteAddr_T_6; // @[Mux.scala 101:16]
  assign GRF_Module_io_WE = io_WEGRF; // @[DataPath.scala 48:22]
  assign GRF_Module_io_WD = _GRFWrite_T ? ALU_Module_io_O : _GRFWrite_T_6; // @[Mux.scala 101:16]
  assign GRF_Module_io_PC = IFU_Module_io_PC; // @[DataPath.scala 50:22]
  assign ALU_Module_io_A1 = GRF_Module_io_O1; // @[DataPath.scala 55:22]
  assign ALU_Module_io_A2 = _ALURead2_T ? GRF_Module_io_O2 : _ALURead2_T_2; // @[Mux.scala 101:16]
  assign ALU_Module_io_ALUOp = io_ALUOp; // @[DataPath.scala 57:25]
  assign DM_Module_clock = clock;
  assign DM_Module_reset = reset;
  assign DM_Module_io_Addr = ALU_Module_io_O; // @[DataPath.scala 59:23]
  assign DM_Module_io_WD = GRF_Module_io_O2; // @[DataPath.scala 60:21]
  assign DM_Module_io_WE = io_WEDM; // @[DataPath.scala 61:21]
  assign DM_Module_io_PC = IFU_Module_io_PC; // @[DataPath.scala 62:21]
  assign EXT_Module_io_imm16 = IFU_Module_io_instr[15:0]; // @[DataPath.scala 64:47]
  assign EXT_Module_io_IsSignEXT = io_IsSignExt; // @[DataPath.scala 65:29]
endmodule
module MIPS(
  input   clock,
  input   reset
);
  wire [31:0] CU_Module_io_instr; // @[MIPS.scala 6:31]
  wire  CU_Module_io_IsEq; // @[MIPS.scala 6:31]
  wire [3:0] CU_Module_io_ALUOp; // @[MIPS.scala 6:31]
  wire  CU_Module_io_WEGRF; // @[MIPS.scala 6:31]
  wire  CU_Module_io_WEDM; // @[MIPS.scala 6:31]
  wire  CU_Module_io_IsBranchType; // @[MIPS.scala 6:31]
  wire  CU_Module_io_IsJType; // @[MIPS.scala 6:31]
  wire  CU_Module_io_IsJr; // @[MIPS.scala 6:31]
  wire  CU_Module_io_ALUSrc; // @[MIPS.scala 6:31]
  wire [1:0] CU_Module_io_WhichToReg; // @[MIPS.scala 6:31]
  wire [1:0] CU_Module_io_RegDst; // @[MIPS.scala 6:31]
  wire  CU_Module_io_IsSignExt; // @[MIPS.scala 6:31]
  wire  DataPath_Module_clock; // @[MIPS.scala 7:43]
  wire  DataPath_Module_reset; // @[MIPS.scala 7:43]
  wire  DataPath_Module_io_WEGRF; // @[MIPS.scala 7:43]
  wire  DataPath_Module_io_WEDM; // @[MIPS.scala 7:43]
  wire [1:0] DataPath_Module_io_RegDst; // @[MIPS.scala 7:43]
  wire [1:0] DataPath_Module_io_WhichToReg; // @[MIPS.scala 7:43]
  wire [3:0] DataPath_Module_io_ALUOp; // @[MIPS.scala 7:43]
  wire  DataPath_Module_io_ALUSrc; // @[MIPS.scala 7:43]
  wire  DataPath_Module_io_IsSignExt; // @[MIPS.scala 7:43]
  wire  DataPath_Module_io_IsBranchType; // @[MIPS.scala 7:43]
  wire  DataPath_Module_io_IsJType; // @[MIPS.scala 7:43]
  wire  DataPath_Module_io_IsJr; // @[MIPS.scala 7:43]
  wire [31:0] DataPath_Module_io_instr; // @[MIPS.scala 7:43]
  wire  DataPath_Module_io_IsEq; // @[MIPS.scala 7:43]
  CU CU_Module ( // @[MIPS.scala 6:31]
    .io_instr(CU_Module_io_instr),
    .io_IsEq(CU_Module_io_IsEq),
    .io_ALUOp(CU_Module_io_ALUOp),
    .io_WEGRF(CU_Module_io_WEGRF),
    .io_WEDM(CU_Module_io_WEDM),
    .io_IsBranchType(CU_Module_io_IsBranchType),
    .io_IsJType(CU_Module_io_IsJType),
    .io_IsJr(CU_Module_io_IsJr),
    .io_ALUSrc(CU_Module_io_ALUSrc),
    .io_WhichToReg(CU_Module_io_WhichToReg),
    .io_RegDst(CU_Module_io_RegDst),
    .io_IsSignExt(CU_Module_io_IsSignExt)
  );
  DataPath DataPath_Module ( // @[MIPS.scala 7:43]
    .clock(DataPath_Module_clock),
    .reset(DataPath_Module_reset),
    .io_WEGRF(DataPath_Module_io_WEGRF),
    .io_WEDM(DataPath_Module_io_WEDM),
    .io_RegDst(DataPath_Module_io_RegDst),
    .io_WhichToReg(DataPath_Module_io_WhichToReg),
    .io_ALUOp(DataPath_Module_io_ALUOp),
    .io_ALUSrc(DataPath_Module_io_ALUSrc),
    .io_IsSignExt(DataPath_Module_io_IsSignExt),
    .io_IsBranchType(DataPath_Module_io_IsBranchType),
    .io_IsJType(DataPath_Module_io_IsJType),
    .io_IsJr(DataPath_Module_io_IsJr),
    .io_instr(DataPath_Module_io_instr),
    .io_IsEq(DataPath_Module_io_IsEq)
  );
  assign CU_Module_io_instr = DataPath_Module_io_instr; // @[MIPS.scala 8:18]
  assign CU_Module_io_IsEq = DataPath_Module_io_IsEq; // @[MIPS.scala 8:18]
  assign DataPath_Module_clock = clock;
  assign DataPath_Module_reset = reset;
  assign DataPath_Module_io_WEGRF = CU_Module_io_WEGRF; // @[MIPS.scala 8:18]
  assign DataPath_Module_io_WEDM = CU_Module_io_WEDM; // @[MIPS.scala 8:18]
  assign DataPath_Module_io_RegDst = CU_Module_io_RegDst; // @[MIPS.scala 8:18]
  assign DataPath_Module_io_WhichToReg = CU_Module_io_WhichToReg; // @[MIPS.scala 8:18]
  assign DataPath_Module_io_ALUOp = CU_Module_io_ALUOp; // @[MIPS.scala 8:18]
  assign DataPath_Module_io_ALUSrc = CU_Module_io_ALUSrc; // @[MIPS.scala 8:18]
  assign DataPath_Module_io_IsSignExt = CU_Module_io_IsSignExt; // @[MIPS.scala 8:18]
  assign DataPath_Module_io_IsBranchType = CU_Module_io_IsBranchType; // @[MIPS.scala 8:18]
  assign DataPath_Module_io_IsJType = CU_Module_io_IsJType; // @[MIPS.scala 8:18]
  assign DataPath_Module_io_IsJr = CU_Module_io_IsJr; // @[MIPS.scala 8:18]
endmodule
